
// Flip-flop.

module smul_flipflop (
    input  wire clk,
    input  wire clken,
    input  wire d,
    output reg  q );

always @(posedge clk)
begin
    if (clken)
        q <= d;
end

endmodule


// Inverter.

module smul_inverter (
    input  wire d,
    output wire q );

assign q = ~d;

endmodule


// Half-adder.

module smul_half_add (
    input  wire x,
    input  wire y,
    output wire d,
    output wire c );

assign d = x ^ y;
assign c = x & y;

endmodule


// Full-adder.

module smul_full_add (
    input  wire x,
    input  wire y,
    input  wire z,
    output wire d,
    output wire c );

assign d = x ^ y ^ z;
assign c = (x & y) | (y & z) | (x & z);

endmodule


// Booth negative flag.

module smul_booth_neg (
    input  wire p0,
    input  wire p1,
    input  wire p2,
    output wire f );

assign f = p2 & ((~p1) | (~p0));

endmodule


// Booth partial product generator.

module smul_booth_prod (
    input  wire p0,
    input  wire p1,
    input  wire p2,
    input  wire u0,
    input  wire u1,
    output reg  y );

always @ (*)
begin
    case ({p2, p1, p0})
        3'b000  : y = 1'b0;
        3'b001  : y = u1;
        3'b010  : y = u1;
        3'b011  : y = u0;
        3'b100  : y = ~u0;
        3'b101  : y = ~u1;
        3'b110  : y = ~u1;
        default : y = 1'b0;
    endcase
end

endmodule


// Deterimine carry generate and carry propagate.

module smul_carry_prop (
    input  wire a,
    input  wire b,
    output wire g,
    output wire p );

assign g = a & b;
assign p = a ^ b;

endmodule


// Merge two carry propagation trees.

module smul_carry_merge (
    input  wire g0,
    input  wire p0,
    input  wire g1,
    input  wire p1,
    output wire g,
    output wire p );

assign g = g1 | (g0 & p1);
assign p = p0 & p1;

endmodule


// Calculate carry-out through a carry propagation tree.

module smul_carry_eval (
    input  wire g,
    input  wire p,
    input  wire cin,
    output wire cout );

assign cout = g | (p & cin);

endmodule

/*
 * 32 x 32 bit fixed point multiplier
 *
 * 0 cycles pipeline delay
 */

module rad4_fixp(
    input  wire [31:0] x,
    input  wire [31:0] y,
    output wire [63:0] p );
    
    wire [63:0] p_temp;
    
    rad4_32bit mult(x,y,p_temp);
    
    assign p = p_temp[41:10];
	
endmodule
/*
 * 32 x 32 bit signed multiplier
 *
 * 0 cycles pipeline delay
 */

module rad4_32bit (
    input  wire [31:0] x,
    input  wire [31:0] y,
    output wire [63:0] p );

wire wadd0d;
wire wadd0c;
wire wboothprod2;
wire wboothneg3;
wire wadd4d;
wire wadd4c;
wire wboothprod6;
wire wcarry7;
wire wcarry8g;
wire wcarry8p;
wire wadd10d;
wire wadd10c;
wire wadd12d;
wire wadd12c;
wire wboothprod14;
wire wboothprod15;
wire wboothneg16;
wire wcarry17;
wire wcarry18g;
wire wcarry18p;
wire wcarry20g;
wire wcarry20p;
wire wadd22d;
wire wadd22c;
wire wadd24d;
wire wadd24c;
wire wboothprod26;
wire wboothprod27;
wire wcarry28;
wire wcarry29g;
wire wcarry29p;
wire wadd31d;
wire wadd31c;
wire wadd33d;
wire wadd33c;
wire wadd35d;
wire wadd35c;
wire wboothprod37;
wire wboothprod38;
wire wboothprod39;
wire wboothneg40;
wire wcarry41;
wire wcarry42g;
wire wcarry42p;
wire wcarry44g;
wire wcarry44p;
wire wcarry46g;
wire wcarry46p;
wire wadd48d;
wire wadd48c;
wire wadd50d;
wire wadd50c;
wire wadd52d;
wire wadd52c;
wire wboothprod54;
wire wboothprod55;
wire wboothprod56;
wire wcarry57;
wire wcarry58g;
wire wcarry58p;
wire wadd60d;
wire wadd60c;
wire wadd62d;
wire wadd62c;
wire wadd64d;
wire wadd64c;
wire wboothprod66;
wire wboothprod67;
wire wboothprod68;
wire wadd69d;
wire wadd69c;
wire wboothprod71;
wire wboothneg72;
wire wcarry73;
wire wcarry74g;
wire wcarry74p;
wire wcarry76g;
wire wcarry76p;
wire wadd78d;
wire wadd78c;
wire wadd80d;
wire wadd80c;
wire wadd82d;
wire wadd82c;
wire wadd84d;
wire wadd84c;
wire wboothprod86;
wire wboothprod87;
wire wboothprod88;
wire wboothprod89;
wire wcarry90;
wire wcarry91g;
wire wcarry91p;
wire wadd93d;
wire wadd93c;
wire wadd95d;
wire wadd95c;
wire wadd97d;
wire wadd97c;
wire wadd99d;
wire wadd99c;
wire wboothprod101;
wire wboothprod102;
wire wboothprod103;
wire wadd104d;
wire wadd104c;
wire wboothprod106;
wire wboothprod107;
wire wboothneg108;
wire wcarry109;
wire wcarry110g;
wire wcarry110p;
wire wcarry112g;
wire wcarry112p;
wire wcarry114g;
wire wcarry114p;
wire wcarry116g;
wire wcarry116p;
wire wadd118d;
wire wadd118c;
wire wadd120d;
wire wadd120c;
wire wadd122d;
wire wadd122c;
wire wadd124d;
wire wadd124c;
wire wboothprod126;
wire wboothprod127;
wire wboothprod128;
wire wadd129d;
wire wadd129c;
wire wboothprod131;
wire wboothprod132;
wire wcarry133;
wire wcarry134g;
wire wcarry134p;
wire wadd136d;
wire wadd136c;
wire wadd138d;
wire wadd138c;
wire wadd140d;
wire wadd140c;
wire wadd142d;
wire wadd142c;
wire wadd144d;
wire wadd144c;
wire wboothprod146;
wire wboothprod147;
wire wboothprod148;
wire wadd149d;
wire wadd149c;
wire wboothprod151;
wire wboothprod152;
wire wboothprod153;
wire wboothneg154;
wire wcarry155;
wire wcarry156g;
wire wcarry156p;
wire wcarry158g;
wire wcarry158p;
wire wadd160d;
wire wadd160c;
wire wadd162d;
wire wadd162c;
wire wadd164d;
wire wadd164c;
wire wadd166d;
wire wadd166c;
wire wadd168d;
wire wadd168c;
wire wboothprod170;
wire wboothprod171;
wire wboothprod172;
wire wadd173d;
wire wadd173c;
wire wboothprod175;
wire wboothprod176;
wire wboothprod177;
wire wcarry178;
wire wcarry179g;
wire wcarry179p;
wire wadd181d;
wire wadd181c;
wire wadd183d;
wire wadd183c;
wire wadd185d;
wire wadd185c;
wire wadd187d;
wire wadd187c;
wire wadd189d;
wire wadd189c;
wire wboothprod191;
wire wboothprod192;
wire wboothprod193;
wire wadd194d;
wire wadd194c;
wire wadd196d;
wire wadd196c;
wire wboothprod198;
wire wboothprod199;
wire wboothprod200;
wire wboothprod201;
wire wboothneg202;
wire wcarry203;
wire wcarry204g;
wire wcarry204p;
wire wcarry206g;
wire wcarry206p;
wire wcarry208g;
wire wcarry208p;
wire wadd210d;
wire wadd210c;
wire wadd212d;
wire wadd212c;
wire wadd214d;
wire wadd214c;
wire wadd216d;
wire wadd216c;
wire wadd218d;
wire wadd218c;
wire wboothprod220;
wire wboothprod221;
wire wboothprod222;
wire wadd223d;
wire wadd223c;
wire wadd225d;
wire wadd225c;
wire wboothprod227;
wire wboothprod228;
wire wboothprod229;
wire wboothprod230;
wire wcarry231;
wire wcarry232g;
wire wcarry232p;
wire wadd234d;
wire wadd234c;
wire wadd236d;
wire wadd236c;
wire wadd238d;
wire wadd238c;
wire wadd240d;
wire wadd240c;
wire wadd242d;
wire wadd242c;
wire wboothprod244;
wire wboothprod245;
wire wboothprod246;
wire wadd247d;
wire wadd247c;
wire wadd249d;
wire wadd249c;
wire wboothprod251;
wire wboothprod252;
wire wboothprod253;
wire wadd254d;
wire wadd254c;
wire wboothprod256;
wire wboothprod257;
wire wboothneg258;
wire wcarry259;
wire wcarry260g;
wire wcarry260p;
wire wcarry262g;
wire wcarry262p;
wire wadd264d;
wire wadd264c;
wire wadd266d;
wire wadd266c;
wire wadd268d;
wire wadd268c;
wire wadd270d;
wire wadd270c;
wire wadd272d;
wire wadd272c;
wire wadd274d;
wire wadd274c;
wire wboothprod276;
wire wboothprod277;
wire wboothprod278;
wire wadd279d;
wire wadd279c;
wire wboothprod281;
wire wboothprod282;
wire wboothprod283;
wire wadd284d;
wire wadd284c;
wire wboothprod286;
wire wboothprod287;
wire wcarry288;
wire wcarry289g;
wire wcarry289p;
wire wadd291d;
wire wadd291c;
wire wadd293d;
wire wadd293c;
wire wadd295d;
wire wadd295c;
wire wadd297d;
wire wadd297c;
wire wadd299d;
wire wadd299c;
wire wadd301d;
wire wadd301c;
wire wadd303d;
wire wadd303c;
wire wboothprod305;
wire wboothprod306;
wire wboothprod307;
wire wadd308d;
wire wadd308c;
wire wboothprod310;
wire wboothprod311;
wire wboothprod312;
wire wadd313d;
wire wadd313c;
wire wboothprod315;
wire wboothprod316;
wire wboothprod317;
wire wboothneg318;
wire wcarry319;
wire wcarry320g;
wire wcarry320p;
wire wcarry322g;
wire wcarry322p;
wire wcarry324g;
wire wcarry324p;
wire wcarry326g;
wire wcarry326p;
wire wcarry328g;
wire wcarry328p;
wire wadd330d;
wire wadd330c;
wire wadd332d;
wire wadd332c;
wire wadd334d;
wire wadd334c;
wire wadd336d;
wire wadd336c;
wire wadd338d;
wire wadd338c;
wire wadd340d;
wire wadd340c;
wire wadd342d;
wire wadd342c;
wire wboothprod344;
wire wboothprod345;
wire wboothprod346;
wire wadd347d;
wire wadd347c;
wire wboothprod349;
wire wboothprod350;
wire wboothprod351;
wire wadd352d;
wire wadd352c;
wire wboothprod354;
wire wboothprod355;
wire wboothprod356;
wire wcarry357;
wire wcarry358g;
wire wcarry358p;
wire wadd360d;
wire wadd360c;
wire wadd362d;
wire wadd362c;
wire wadd364d;
wire wadd364c;
wire wadd366d;
wire wadd366c;
wire wadd368d;
wire wadd368c;
wire wadd370d;
wire wadd370c;
wire wadd372d;
wire wadd372c;
wire wadd374d;
wire wadd374c;
wire wboothprod376;
wire wboothprod377;
wire wboothprod378;
wire wadd379d;
wire wadd379c;
wire wboothprod381;
wire wboothprod382;
wire wboothprod383;
wire wadd384d;
wire wadd384c;
wire wboothprod386;
wire wboothprod387;
wire wboothprod388;
wire wboothprod389;
wire wboothneg390;
wire wcarry391;
wire wcarry392g;
wire wcarry392p;
wire wcarry394g;
wire wcarry394p;
wire wadd396d;
wire wadd396c;
wire wadd398d;
wire wadd398c;
wire wadd400d;
wire wadd400c;
wire wadd402d;
wire wadd402c;
wire wadd404d;
wire wadd404c;
wire wadd406d;
wire wadd406c;
wire wadd408d;
wire wadd408c;
wire wadd410d;
wire wadd410c;
wire wboothprod412;
wire wboothprod413;
wire wboothprod414;
wire wadd415d;
wire wadd415c;
wire wboothprod417;
wire wboothprod418;
wire wboothprod419;
wire wadd420d;
wire wadd420c;
wire wboothprod422;
wire wboothprod423;
wire wboothprod424;
wire wboothprod425;
wire wcarry426;
wire wcarry427g;
wire wcarry427p;
wire wadd429d;
wire wadd429c;
wire wadd431d;
wire wadd431c;
wire wadd433d;
wire wadd433c;
wire wadd435d;
wire wadd435c;
wire wadd437d;
wire wadd437c;
wire wadd439d;
wire wadd439c;
wire wadd441d;
wire wadd441c;
wire wadd443d;
wire wadd443c;
wire wboothprod445;
wire wboothprod446;
wire wboothprod447;
wire wadd448d;
wire wadd448c;
wire wboothprod450;
wire wboothprod451;
wire wboothprod452;
wire wadd453d;
wire wadd453c;
wire wboothprod455;
wire wboothprod456;
wire wboothprod457;
wire wadd458d;
wire wadd458c;
wire wboothprod460;
wire wboothprod461;
wire wboothneg462;
wire wcarry463;
wire wcarry464g;
wire wcarry464p;
wire wcarry466g;
wire wcarry466p;
wire wcarry468g;
wire wcarry468p;
wire wadd470d;
wire wadd470c;
wire wadd472d;
wire wadd472c;
wire wadd474d;
wire wadd474c;
wire wadd476d;
wire wadd476c;
wire wadd478d;
wire wadd478c;
wire wadd480d;
wire wadd480c;
wire wadd482d;
wire wadd482c;
wire wadd484d;
wire wadd484c;
wire wboothprod486;
wire wboothprod487;
wire wboothprod488;
wire wadd489d;
wire wadd489c;
wire wboothprod491;
wire wboothprod492;
wire wboothprod493;
wire wadd494d;
wire wadd494c;
wire wadd496d;
wire wadd496c;
wire wboothprod498;
wire wboothprod499;
wire wboothprod500;
wire wboothprod501;
wire wboothprod502;
wire wcarry503;
wire wcarry504g;
wire wcarry504p;
wire wadd506d;
wire wadd506c;
wire wadd508d;
wire wadd508c;
wire wadd510d;
wire wadd510c;
wire wadd512d;
wire wadd512c;
wire wadd514d;
wire wadd514c;
wire wadd516d;
wire wadd516c;
wire wadd518d;
wire wadd518c;
wire wadd520d;
wire wadd520c;
wire wboothprod522;
wire wboothprod523;
wire wboothprod524;
wire wadd525d;
wire wadd525c;
wire wboothprod527;
wire wboothprod528;
wire wboothprod529;
wire wadd530d;
wire wadd530c;
wire wboothprod532;
wire wboothprod533;
wire wboothprod534;
wire wadd535d;
wire wadd535c;
wire wadd537d;
wire wadd537c;
wire wboothprod539;
wire wboothprod540;
wire wboothprod541;
wire wboothneg542;
wire wcarry543;
wire wcarry544g;
wire wcarry544p;
wire wcarry546g;
wire wcarry546p;
wire wadd548d;
wire wadd548c;
wire wadd550d;
wire wadd550c;
wire wadd552d;
wire wadd552c;
wire wadd554d;
wire wadd554c;
wire wadd556d;
wire wadd556c;
wire wadd558d;
wire wadd558c;
wire wadd560d;
wire wadd560c;
wire wadd562d;
wire wadd562c;
wire wboothprod564;
wire wboothprod565;
wire wboothprod566;
wire wadd567d;
wire wadd567c;
wire wboothprod569;
wire wboothprod570;
wire wboothprod571;
wire wadd572d;
wire wadd572c;
wire wadd574d;
wire wadd574c;
wire wboothprod576;
wire wboothprod577;
wire wboothprod578;
wire wadd579d;
wire wadd579c;
wire wboothprod581;
wire wboothprod582;
wire wboothprod583;
wire wcarry584;
wire wcarry585g;
wire wcarry585p;
wire wadd587d;
wire wadd587c;
wire wadd589d;
wire wadd589c;
wire wadd591d;
wire wadd591c;
wire wadd593d;
wire wadd593c;
wire wadd595d;
wire wadd595c;
wire wadd597d;
wire wadd597c;
wire wadd599d;
wire wadd599c;
wire wadd601d;
wire wadd601c;
wire wboothprod603;
wire wboothprod604;
wire wboothprod605;
wire wadd606d;
wire wadd606c;
wire wboothprod608;
wire wboothprod609;
wire wboothprod610;
wire wadd611d;
wire wadd611c;
wire wadd613d;
wire wadd613c;
wire wboothprod615;
wire wboothprod616;
wire wboothprod617;
wire wadd618d;
wire wadd618c;
wire wboothprod620;
wire wboothprod621;
wire wboothprod622;
wire wadd623d;
wire wadd623c;
wire wboothprod625;
wire wboothneg626;
wire wcarry627;
wire wcarry628g;
wire wcarry628p;
wire wcarry630g;
wire wcarry630p;
wire wcarry632g;
wire wcarry632p;
wire wcarry634g;
wire wcarry634p;
wire wadd636d;
wire wadd636c;
wire wadd638d;
wire wadd638c;
wire wadd640d;
wire wadd640c;
wire wadd642d;
wire wadd642c;
wire wadd644d;
wire wadd644c;
wire wadd646d;
wire wadd646c;
wire wadd648d;
wire wadd648c;
wire wadd650d;
wire wadd650c;
wire wadd652d;
wire wadd652c;
wire wboothprod654;
wire wboothprod655;
wire wboothprod656;
wire wadd657d;
wire wadd657c;
wire wadd659d;
wire wadd659c;
wire wboothprod661;
wire wboothprod662;
wire wboothprod663;
wire wadd664d;
wire wadd664c;
wire wboothprod666;
wire wboothprod667;
wire wboothprod668;
wire wadd669d;
wire wadd669c;
wire wboothprod671;
wire wboothprod672;
wire wboothprod673;
wire wboothprod674;
wire wcarry675;
wire wcarry676g;
wire wcarry676p;
wire wadd678d;
wire wadd678c;
wire wadd680d;
wire wadd680c;
wire wadd682d;
wire wadd682c;
wire wadd684d;
wire wadd684c;
wire wadd686d;
wire wadd686c;
wire wadd688d;
wire wadd688c;
wire wadd690d;
wire wadd690c;
wire wadd692d;
wire wadd692c;
wire wadd694d;
wire wadd694c;
wire wboothprod696;
wire wboothprod697;
wire wboothprod698;
wire wadd699d;
wire wadd699c;
wire wboothprod701;
wire wboothprod702;
wire wboothprod703;
wire wadd704d;
wire wadd704c;
wire wadd706d;
wire wadd706c;
wire wboothprod708;
wire wboothprod709;
wire wboothprod710;
wire wadd711d;
wire wadd711c;
wire wboothprod713;
wire wboothprod714;
wire wboothprod715;
wire wadd716d;
wire wadd716c;
wire wboothprod718;
wire wboothprod719;
wire wboothneg720;
wire wcarry721;
wire wcarry722g;
wire wcarry722p;
wire wcarry724g;
wire wcarry724p;
wire wadd726d;
wire wadd726c;
wire wadd728d;
wire wadd728c;
wire wadd730d;
wire wadd730c;
wire wadd732d;
wire wadd732c;
wire wadd734d;
wire wadd734c;
wire wadd736d;
wire wadd736c;
wire wadd738d;
wire wadd738c;
wire wadd740d;
wire wadd740c;
wire wadd742d;
wire wadd742c;
wire wadd744d;
wire wadd744c;
wire wboothprod746;
wire wboothprod747;
wire wboothprod748;
wire wadd749d;
wire wadd749c;
wire wadd751d;
wire wadd751c;
wire wboothprod753;
wire wboothprod754;
wire wboothprod755;
wire wadd756d;
wire wadd756c;
wire wboothprod758;
wire wboothprod759;
wire wboothprod760;
wire wadd761d;
wire wadd761c;
wire wboothprod763;
wire wboothprod764;
wire wboothprod765;
wire wboothprod766;
wire wboothprod767;
wire wcarry768;
wire wcarry769g;
wire wcarry769p;
wire wadd771d;
wire wadd771c;
wire wadd773d;
wire wadd773c;
wire wadd775d;
wire wadd775c;
wire wadd777d;
wire wadd777c;
wire wadd779d;
wire wadd779c;
wire wadd781d;
wire wadd781c;
wire wadd783d;
wire wadd783c;
wire wadd785d;
wire wadd785c;
wire wadd787d;
wire wadd787c;
wire wadd789d;
wire wadd789c;
wire wboothprod791;
wire wboothprod792;
wire wboothprod793;
wire wadd794d;
wire wadd794c;
wire wboothprod796;
wire wboothprod797;
wire wboothprod798;
wire wadd799d;
wire wadd799c;
wire wadd801d;
wire wadd801c;
wire wboothprod803;
wire wboothprod804;
wire wboothprod805;
wire wadd806d;
wire wadd806c;
wire wboothprod808;
wire wboothprod809;
wire wboothprod810;
wire wadd811d;
wire wadd811c;
wire wboothprod813;
wire wboothprod814;
wire wboothprod815;
wire wboothneg816;
wire wcarry817;
wire wcarry818g;
wire wcarry818p;
wire wcarry820g;
wire wcarry820p;
wire wcarry822g;
wire wcarry822p;
wire wadd824d;
wire wadd824c;
wire wadd826d;
wire wadd826c;
wire wadd828d;
wire wadd828c;
wire wadd830d;
wire wadd830c;
wire wadd832d;
wire wadd832c;
wire wadd834d;
wire wadd834c;
wire wadd836d;
wire wadd836c;
wire wadd838d;
wire wadd838c;
wire wadd840d;
wire wadd840c;
wire wadd842d;
wire wadd842c;
wire wboothprod844;
wire wboothprod845;
wire wboothprod846;
wire wadd847d;
wire wadd847c;
wire wadd849d;
wire wadd849c;
wire wboothprod851;
wire wboothprod852;
wire wboothprod853;
wire wadd854d;
wire wadd854c;
wire wboothprod856;
wire wboothprod857;
wire wboothprod858;
wire wadd859d;
wire wadd859c;
wire wboothprod861;
wire wboothprod862;
wire wboothprod863;
wire wadd864d;
wire wadd864c;
wire wboothprod866;
wire wboothprod867;
wire wboothprod868;
wire wcarry869;
wire wcarry870g;
wire wcarry870p;
wire wadd872d;
wire wadd872c;
wire wadd874d;
wire wadd874c;
wire wadd876d;
wire wadd876c;
wire wadd878d;
wire wadd878c;
wire wadd880d;
wire wadd880c;
wire wadd882d;
wire wadd882c;
wire wadd884d;
wire wadd884c;
wire wadd886d;
wire wadd886c;
wire wadd888d;
wire wadd888c;
wire wadd890d;
wire wadd890c;
wire wboothprod892;
wire wboothprod893;
wire wboothprod894;
wire wadd895d;
wire wadd895c;
wire wadd897d;
wire wadd897c;
wire wboothprod899;
wire wboothprod900;
wire wboothprod901;
wire wadd902d;
wire wadd902c;
wire wboothprod904;
wire wboothprod905;
wire wboothprod906;
wire wadd907d;
wire wadd907c;
wire wboothprod909;
wire wboothprod910;
wire wboothprod911;
wire wadd912d;
wire wadd912c;
wire wadd914d;
wire wadd914c;
wire wboothprod916;
wire wboothprod917;
wire wboothprod918;
wire wboothprod919;
wire wboothneg920;
wire wcarry921;
wire wcarry922g;
wire wcarry922p;
wire wcarry924g;
wire wcarry924p;
wire wadd926d;
wire wadd926c;
wire wadd928d;
wire wadd928c;
wire wadd930d;
wire wadd930c;
wire wadd932d;
wire wadd932c;
wire wadd934d;
wire wadd934c;
wire wadd936d;
wire wadd936c;
wire wadd938d;
wire wadd938c;
wire wadd940d;
wire wadd940c;
wire wadd942d;
wire wadd942c;
wire wadd944d;
wire wadd944c;
wire wboothprod946;
wire wboothprod947;
wire wboothprod948;
wire wadd949d;
wire wadd949c;
wire wadd951d;
wire wadd951c;
wire wadd953d;
wire wadd953c;
wire wboothprod955;
wire wboothprod956;
wire wboothprod957;
wire wadd958d;
wire wadd958c;
wire wboothprod960;
wire wboothprod961;
wire wboothprod962;
wire wadd963d;
wire wadd963c;
wire wboothprod965;
wire wboothprod966;
wire wboothprod967;
wire wadd968d;
wire wadd968c;
wire wboothprod970;
wire wboothprod971;
wire wboothprod972;
wire wboothprod973;
wire wcarry974;
wire wcarry975g;
wire wcarry975p;
wire wadd977d;
wire wadd977c;
wire wadd979d;
wire wadd979c;
wire wadd981d;
wire wadd981c;
wire wadd983d;
wire wadd983c;
wire wadd985d;
wire wadd985c;
wire wadd987d;
wire wadd987c;
wire wadd989d;
wire wadd989c;
wire wadd991d;
wire wadd991c;
wire wadd993d;
wire wadd993c;
wire wadd995d;
wire wadd995c;
wire wboothprod997;
wire wboothprod998;
wire wboothprod999;
wire wadd1000d;
wire wadd1000c;
wire wadd1002d;
wire wadd1002c;
wire wboothprod1004;
wire wboothprod1005;
wire wboothprod1006;
wire wadd1007d;
wire wadd1007c;
wire wboothprod1009;
wire wboothprod1010;
wire wboothprod1011;
wire wadd1012d;
wire wadd1012c;
wire wboothprod1014;
wire wboothprod1015;
wire wboothprod1016;
wire wadd1017d;
wire wadd1017c;
wire wadd1019d;
wire wadd1019c;
wire wboothprod1021;
wire wboothprod1022;
wire wboothprod1023;
wire wboothprod1024;
wire wcarry1025;
wire wcarry1026g;
wire wcarry1026p;
wire wcarry1028g;
wire wcarry1028p;
wire wcarry1030g;
wire wcarry1030p;
wire wcarry1032g;
wire wcarry1032p;
wire wcarry1034g;
wire wcarry1034p;
wire wcarry1036g;
wire wcarry1036p;
wire wadd1038d;
wire wadd1038c;
wire wadd1040d;
wire wadd1040c;
wire wadd1042d;
wire wadd1042c;
wire wadd1044d;
wire wadd1044c;
wire wadd1046d;
wire wadd1046c;
wire wadd1048d;
wire wadd1048c;
wire wadd1050d;
wire wadd1050c;
wire wadd1052d;
wire wadd1052c;
wire wadd1054d;
wire wadd1054c;
wire wadd1056d;
wire wadd1056c;
wire wboothprod1058;
wire wboothprod1059;
wire wadd1060d;
wire wadd1060c;
wire wadd1062d;
wire wadd1062c;
wire wboothprod1064;
wire wboothprod1065;
wire wboothprod1066;
wire wadd1067d;
wire wadd1067c;
wire wboothprod1069;
wire wboothprod1070;
wire wboothprod1071;
wire wadd1072d;
wire wadd1072c;
wire wboothprod1074;
wire wboothprod1075;
wire wboothprod1076;
wire wadd1077d;
wire wadd1077c;
wire wadd1079d;
wire wadd1079c;
wire wboothprod1081;
wire wboothprod1082;
wire wboothprod1083;
wire wboothprod1084;
wire wcarry1085;
wire wcarry1086g;
wire wcarry1086p;
wire wadd1088d;
wire wadd1088c;
wire wadd1090d;
wire wadd1090c;
wire wadd1092d;
wire wadd1092c;
wire wadd1094d;
wire wadd1094c;
wire wadd1096d;
wire wadd1096c;
wire wadd1098d;
wire wadd1098c;
wire wadd1100d;
wire wadd1100c;
wire wadd1102d;
wire wadd1102c;
wire wadd1104d;
wire wadd1104c;
wire wadd1106d;
wire wadd1106c;
wire winv1108;
wire winv1109;
wire wboothprod1110;
wire wboothprod1111;
wire wadd1112d;
wire wadd1112c;
wire wadd1114d;
wire wadd1114c;
wire wboothprod1116;
wire wboothprod1117;
wire wboothprod1118;
wire wadd1119d;
wire wadd1119c;
wire wboothprod1121;
wire wboothprod1122;
wire wboothprod1123;
wire wadd1124d;
wire wadd1124c;
wire wboothprod1126;
wire wboothprod1127;
wire wboothprod1128;
wire wadd1129d;
wire wadd1129c;
wire wadd1131d;
wire wadd1131c;
wire wboothprod1133;
wire wboothprod1134;
wire wboothprod1135;
wire wboothprod1136;
wire wcarry1137;
wire wcarry1138g;
wire wcarry1138p;
wire wcarry1140g;
wire wcarry1140p;
wire wadd1142d;
wire wadd1142c;
wire wadd1144d;
wire wadd1144c;
wire wadd1146d;
wire wadd1146c;
wire wadd1148d;
wire wadd1148c;
wire wadd1150d;
wire wadd1150c;
wire wadd1152d;
wire wadd1152c;
wire wadd1154d;
wire wadd1154c;
wire wadd1156d;
wire wadd1156c;
wire wadd1158d;
wire wadd1158c;
wire wadd1160d;
wire wadd1160c;
wire wboothprod1162;
wire wboothprod1163;
wire wadd1164d;
wire wadd1164c;
wire wadd1166d;
wire wadd1166c;
wire wboothprod1168;
wire wboothprod1169;
wire wboothprod1170;
wire wadd1171d;
wire wadd1171c;
wire wboothprod1173;
wire wboothprod1174;
wire wboothprod1175;
wire wadd1176d;
wire wadd1176c;
wire wboothprod1178;
wire wboothprod1179;
wire wboothprod1180;
wire wadd1181d;
wire wadd1181c;
wire wboothprod1183;
wire wboothprod1184;
wire wboothprod1185;
wire wcarry1186;
wire wcarry1187g;
wire wcarry1187p;
wire wadd1189d;
wire wadd1189c;
wire wadd1191d;
wire wadd1191c;
wire wadd1193d;
wire wadd1193c;
wire wadd1195d;
wire wadd1195c;
wire wadd1197d;
wire wadd1197c;
wire wadd1199d;
wire wadd1199c;
wire wadd1201d;
wire wadd1201c;
wire wadd1203d;
wire wadd1203c;
wire wadd1205d;
wire wadd1205c;
wire wadd1207d;
wire wadd1207c;
wire winv1209;
wire wboothprod1210;
wire wboothprod1211;
wire wboothprod1212;
wire wadd1213d;
wire wadd1213c;
wire wadd1215d;
wire wadd1215c;
wire wboothprod1217;
wire wboothprod1218;
wire wboothprod1219;
wire wadd1220d;
wire wadd1220c;
wire wboothprod1222;
wire wboothprod1223;
wire wboothprod1224;
wire wadd1225d;
wire wadd1225c;
wire wboothprod1227;
wire wboothprod1228;
wire wboothprod1229;
wire wboothprod1230;
wire wboothprod1231;
wire wcarry1232;
wire wcarry1233g;
wire wcarry1233p;
wire wcarry1235g;
wire wcarry1235p;
wire wcarry1237g;
wire wcarry1237p;
wire wadd1239d;
wire wadd1239c;
wire wadd1241d;
wire wadd1241c;
wire wadd1243d;
wire wadd1243c;
wire wadd1245d;
wire wadd1245c;
wire wadd1247d;
wire wadd1247c;
wire wadd1249d;
wire wadd1249c;
wire wadd1251d;
wire wadd1251c;
wire wadd1253d;
wire wadd1253c;
wire wadd1255d;
wire wadd1255c;
wire wboothprod1257;
wire wboothprod1258;
wire wadd1259d;
wire wadd1259c;
wire wboothprod1261;
wire wboothprod1262;
wire wboothprod1263;
wire wadd1264d;
wire wadd1264c;
wire wadd1266d;
wire wadd1266c;
wire wboothprod1268;
wire wboothprod1269;
wire wboothprod1270;
wire wadd1271d;
wire wadd1271c;
wire wboothprod1273;
wire wboothprod1274;
wire wboothprod1275;
wire wadd1276d;
wire wadd1276c;
wire wboothprod1278;
wire wboothprod1279;
wire wcarry1280;
wire wcarry1281g;
wire wcarry1281p;
wire wadd1283d;
wire wadd1283c;
wire wadd1285d;
wire wadd1285c;
wire wadd1287d;
wire wadd1287c;
wire wadd1289d;
wire wadd1289c;
wire wadd1291d;
wire wadd1291c;
wire wadd1293d;
wire wadd1293c;
wire wadd1295d;
wire wadd1295c;
wire wadd1297d;
wire wadd1297c;
wire wadd1299d;
wire wadd1299c;
wire wadd1301d;
wire wadd1301c;
wire winv1303;
wire wboothprod1304;
wire wboothprod1305;
wire wboothprod1306;
wire wadd1307d;
wire wadd1307c;
wire wadd1309d;
wire wadd1309c;
wire wboothprod1311;
wire wboothprod1312;
wire wboothprod1313;
wire wadd1314d;
wire wadd1314c;
wire wboothprod1316;
wire wboothprod1317;
wire wboothprod1318;
wire wadd1319d;
wire wadd1319c;
wire wboothprod1321;
wire wboothprod1322;
wire wboothprod1323;
wire wboothprod1324;
wire wcarry1325;
wire wcarry1326g;
wire wcarry1326p;
wire wcarry1328g;
wire wcarry1328p;
wire wadd1330d;
wire wadd1330c;
wire wadd1332d;
wire wadd1332c;
wire wadd1334d;
wire wadd1334c;
wire wadd1336d;
wire wadd1336c;
wire wadd1338d;
wire wadd1338c;
wire wadd1340d;
wire wadd1340c;
wire wadd1342d;
wire wadd1342c;
wire wadd1344d;
wire wadd1344c;
wire wadd1346d;
wire wadd1346c;
wire wboothprod1348;
wire wboothprod1349;
wire wadd1350d;
wire wadd1350c;
wire wboothprod1352;
wire wboothprod1353;
wire wboothprod1354;
wire wadd1355d;
wire wadd1355c;
wire wadd1357d;
wire wadd1357c;
wire wboothprod1359;
wire wboothprod1360;
wire wboothprod1361;
wire wadd1362d;
wire wadd1362c;
wire wboothprod1364;
wire wboothprod1365;
wire wboothprod1366;
wire wboothprod1367;
wire wcarry1368;
wire wcarry1369g;
wire wcarry1369p;
wire wadd1371d;
wire wadd1371c;
wire wadd1373d;
wire wadd1373c;
wire wadd1375d;
wire wadd1375c;
wire wadd1377d;
wire wadd1377c;
wire wadd1379d;
wire wadd1379c;
wire wadd1381d;
wire wadd1381c;
wire wadd1383d;
wire wadd1383c;
wire wadd1385d;
wire wadd1385c;
wire wadd1387d;
wire wadd1387c;
wire winv1389;
wire wboothprod1390;
wire wboothprod1391;
wire wboothprod1392;
wire wadd1393d;
wire wadd1393c;
wire wboothprod1395;
wire wboothprod1396;
wire wboothprod1397;
wire wadd1398d;
wire wadd1398c;
wire wadd1400d;
wire wadd1400c;
wire wboothprod1402;
wire wboothprod1403;
wire wboothprod1404;
wire wadd1405d;
wire wadd1405c;
wire wboothprod1407;
wire wboothprod1408;
wire wboothprod1409;
wire wcarry1410;
wire wcarry1411g;
wire wcarry1411p;
wire wcarry1413g;
wire wcarry1413p;
wire wcarry1415g;
wire wcarry1415p;
wire wcarry1417g;
wire wcarry1417p;
wire wadd1419d;
wire wadd1419c;
wire wadd1421d;
wire wadd1421c;
wire wadd1423d;
wire wadd1423c;
wire wadd1425d;
wire wadd1425c;
wire wadd1427d;
wire wadd1427c;
wire wadd1429d;
wire wadd1429c;
wire wadd1431d;
wire wadd1431c;
wire wadd1433d;
wire wadd1433c;
wire wadd1435d;
wire wadd1435c;
wire wboothprod1437;
wire wboothprod1438;
wire wadd1439d;
wire wadd1439c;
wire wboothprod1441;
wire wboothprod1442;
wire wboothprod1443;
wire wadd1444d;
wire wadd1444c;
wire wadd1446d;
wire wadd1446c;
wire wboothprod1448;
wire wboothprod1449;
wire wboothprod1450;
wire wadd1451d;
wire wadd1451c;
wire wboothprod1453;
wire wboothprod1454;
wire wboothprod1455;
wire wcarry1456;
wire wcarry1457g;
wire wcarry1457p;
wire wadd1459d;
wire wadd1459c;
wire wadd1461d;
wire wadd1461c;
wire wadd1463d;
wire wadd1463c;
wire wadd1465d;
wire wadd1465c;
wire wadd1467d;
wire wadd1467c;
wire wadd1469d;
wire wadd1469c;
wire wadd1471d;
wire wadd1471c;
wire wadd1473d;
wire wadd1473c;
wire wadd1475d;
wire wadd1475c;
wire winv1477;
wire wboothprod1478;
wire wboothprod1479;
wire wboothprod1480;
wire wadd1481d;
wire wadd1481c;
wire wboothprod1483;
wire wboothprod1484;
wire wboothprod1485;
wire wadd1486d;
wire wadd1486c;
wire wadd1488d;
wire wadd1488c;
wire wboothprod1490;
wire wboothprod1491;
wire wboothprod1492;
wire wboothprod1493;
wire wboothprod1494;
wire wcarry1495;
wire wcarry1496g;
wire wcarry1496p;
wire wcarry1498g;
wire wcarry1498p;
wire wadd1500d;
wire wadd1500c;
wire wadd1502d;
wire wadd1502c;
wire wadd1504d;
wire wadd1504c;
wire wadd1506d;
wire wadd1506c;
wire wadd1508d;
wire wadd1508c;
wire wadd1510d;
wire wadd1510c;
wire wadd1512d;
wire wadd1512c;
wire wadd1514d;
wire wadd1514c;
wire wadd1516d;
wire wadd1516c;
wire wboothprod1518;
wire wboothprod1519;
wire wadd1520d;
wire wadd1520c;
wire wboothprod1522;
wire wboothprod1523;
wire wboothprod1524;
wire wadd1525d;
wire wadd1525c;
wire wboothprod1527;
wire wboothprod1528;
wire wboothprod1529;
wire wadd1530d;
wire wadd1530c;
wire wboothprod1532;
wire wboothprod1533;
wire wcarry1534;
wire wcarry1535g;
wire wcarry1535p;
wire wadd1537d;
wire wadd1537c;
wire wadd1539d;
wire wadd1539c;
wire wadd1541d;
wire wadd1541c;
wire wadd1543d;
wire wadd1543c;
wire wadd1545d;
wire wadd1545c;
wire wadd1547d;
wire wadd1547c;
wire wadd1549d;
wire wadd1549c;
wire wadd1551d;
wire wadd1551c;
wire wadd1553d;
wire wadd1553c;
wire winv1555;
wire wboothprod1556;
wire wboothprod1557;
wire wboothprod1558;
wire wadd1559d;
wire wadd1559c;
wire wboothprod1561;
wire wboothprod1562;
wire wboothprod1563;
wire wadd1564d;
wire wadd1564c;
wire wboothprod1566;
wire wboothprod1567;
wire wboothprod1568;
wire wboothprod1569;
wire wcarry1570;
wire wcarry1571g;
wire wcarry1571p;
wire wcarry1573g;
wire wcarry1573p;
wire wcarry1575g;
wire wcarry1575p;
wire wadd1577d;
wire wadd1577c;
wire wadd1579d;
wire wadd1579c;
wire wadd1581d;
wire wadd1581c;
wire wadd1583d;
wire wadd1583c;
wire wadd1585d;
wire wadd1585c;
wire wadd1587d;
wire wadd1587c;
wire wadd1589d;
wire wadd1589c;
wire wadd1591d;
wire wadd1591c;
wire wadd1593d;
wire wadd1593c;
wire wboothprod1595;
wire wboothprod1596;
wire wadd1597d;
wire wadd1597c;
wire wboothprod1599;
wire wboothprod1600;
wire wboothprod1601;
wire wadd1602d;
wire wadd1602c;
wire wboothprod1604;
wire wboothprod1605;
wire wboothprod1606;
wire wboothprod1607;
wire wcarry1608;
wire wcarry1609g;
wire wcarry1609p;
wire wadd1611d;
wire wadd1611c;
wire wadd1613d;
wire wadd1613c;
wire wadd1615d;
wire wadd1615c;
wire wadd1617d;
wire wadd1617c;
wire wadd1619d;
wire wadd1619c;
wire wadd1621d;
wire wadd1621c;
wire wadd1623d;
wire wadd1623c;
wire wadd1625d;
wire wadd1625c;
wire winv1627;
wire wboothprod1628;
wire wboothprod1629;
wire wboothprod1630;
wire wadd1631d;
wire wadd1631c;
wire wboothprod1633;
wire wboothprod1634;
wire wboothprod1635;
wire wadd1636d;
wire wadd1636c;
wire wboothprod1638;
wire wboothprod1639;
wire wboothprod1640;
wire wcarry1641;
wire wcarry1642g;
wire wcarry1642p;
wire wcarry1644g;
wire wcarry1644p;
wire wadd1646d;
wire wadd1646c;
wire wadd1648d;
wire wadd1648c;
wire wadd1650d;
wire wadd1650c;
wire wadd1652d;
wire wadd1652c;
wire wadd1654d;
wire wadd1654c;
wire wadd1656d;
wire wadd1656c;
wire wadd1658d;
wire wadd1658c;
wire wboothprod1660;
wire wboothprod1661;
wire wadd1662d;
wire wadd1662c;
wire wboothprod1664;
wire wboothprod1665;
wire wboothprod1666;
wire wadd1667d;
wire wadd1667c;
wire wboothprod1669;
wire wboothprod1670;
wire wboothprod1671;
wire wcarry1672;
wire wcarry1673g;
wire wcarry1673p;
wire wadd1675d;
wire wadd1675c;
wire wadd1677d;
wire wadd1677c;
wire wadd1679d;
wire wadd1679c;
wire wadd1681d;
wire wadd1681c;
wire wadd1683d;
wire wadd1683c;
wire wadd1685d;
wire wadd1685c;
wire wadd1687d;
wire wadd1687c;
wire winv1689;
wire wboothprod1690;
wire wboothprod1691;
wire wboothprod1692;
wire wadd1693d;
wire wadd1693c;
wire wboothprod1695;
wire wboothprod1696;
wire wboothprod1697;
wire wadd1698d;
wire wadd1698c;
wire wboothprod1700;
wire wboothprod1701;
wire wcarry1702;
wire wcarry1703g;
wire wcarry1703p;
wire wcarry1705g;
wire wcarry1705p;
wire wcarry1707g;
wire wcarry1707p;
wire wcarry1709g;
wire wcarry1709p;
wire wcarry1711g;
wire wcarry1711p;
wire wadd1713d;
wire wadd1713c;
wire wadd1715d;
wire wadd1715c;
wire wadd1717d;
wire wadd1717c;
wire wadd1719d;
wire wadd1719c;
wire wadd1721d;
wire wadd1721c;
wire wadd1723d;
wire wadd1723c;
wire wadd1725d;
wire wadd1725c;
wire wboothprod1727;
wire wboothprod1728;
wire wadd1729d;
wire wadd1729c;
wire wboothprod1731;
wire wboothprod1732;
wire wboothprod1733;
wire wadd1734d;
wire wadd1734c;
wire wboothprod1736;
wire wboothprod1737;
wire wcarry1738;
wire wcarry1739g;
wire wcarry1739p;
wire wadd1741d;
wire wadd1741c;
wire wadd1743d;
wire wadd1743c;
wire wadd1745d;
wire wadd1745c;
wire wadd1747d;
wire wadd1747c;
wire wadd1749d;
wire wadd1749c;
wire wadd1751d;
wire wadd1751c;
wire wadd1753d;
wire wadd1753c;
wire winv1755;
wire wboothprod1756;
wire wboothprod1757;
wire wboothprod1758;
wire wadd1759d;
wire wadd1759c;
wire wboothprod1761;
wire wboothprod1762;
wire wboothprod1763;
wire wboothprod1764;
wire wcarry1765;
wire wcarry1766g;
wire wcarry1766p;
wire wcarry1768g;
wire wcarry1768p;
wire wadd1770d;
wire wadd1770c;
wire wadd1772d;
wire wadd1772c;
wire wadd1774d;
wire wadd1774c;
wire wadd1776d;
wire wadd1776c;
wire wadd1778d;
wire wadd1778c;
wire wadd1780d;
wire wadd1780c;
wire wboothprod1782;
wire wboothprod1783;
wire wadd1784d;
wire wadd1784c;
wire wadd1786d;
wire wadd1786c;
wire wboothprod1788;
wire wboothprod1789;
wire wboothprod1790;
wire wboothprod1791;
wire wcarry1792;
wire wcarry1793g;
wire wcarry1793p;
wire wadd1795d;
wire wadd1795c;
wire wadd1797d;
wire wadd1797c;
wire wadd1799d;
wire wadd1799c;
wire wadd1801d;
wire wadd1801c;
wire wadd1803d;
wire wadd1803c;
wire wadd1805d;
wire wadd1805c;
wire winv1807;
wire wboothprod1808;
wire wboothprod1809;
wire wboothprod1810;
wire wadd1811d;
wire wadd1811c;
wire wboothprod1813;
wire wboothprod1814;
wire wboothprod1815;
wire wcarry1816;
wire wcarry1817g;
wire wcarry1817p;
wire wcarry1819g;
wire wcarry1819p;
wire wcarry1821g;
wire wcarry1821p;
wire wadd1823d;
wire wadd1823c;
wire wadd1825d;
wire wadd1825c;
wire wadd1827d;
wire wadd1827c;
wire wadd1829d;
wire wadd1829c;
wire wadd1831d;
wire wadd1831c;
wire wboothprod1833;
wire wboothprod1834;
wire wadd1835d;
wire wadd1835c;
wire wboothprod1837;
wire wboothprod1838;
wire wboothprod1839;
wire wcarry1840;
wire wcarry1841g;
wire wcarry1841p;
wire wadd1843d;
wire wadd1843c;
wire wadd1845d;
wire wadd1845c;
wire wadd1847d;
wire wadd1847c;
wire wadd1849d;
wire wadd1849c;
wire wadd1851d;
wire wadd1851c;
wire winv1853;
wire wboothprod1854;
wire wboothprod1855;
wire wboothprod1856;
wire wadd1857d;
wire wadd1857c;
wire wboothprod1859;
wire wboothprod1860;
wire wcarry1861;
wire wcarry1862g;
wire wcarry1862p;
wire wcarry1864g;
wire wcarry1864p;
wire wadd1866d;
wire wadd1866c;
wire wadd1868d;
wire wadd1868c;
wire wadd1870d;
wire wadd1870c;
wire wadd1872d;
wire wadd1872c;
wire wadd1874d;
wire wadd1874c;
wire wboothprod1876;
wire wboothprod1877;
wire wadd1878d;
wire wadd1878c;
wire wboothprod1880;
wire wboothprod1881;
wire wcarry1882;
wire wcarry1883g;
wire wcarry1883p;
wire wadd1885d;
wire wadd1885c;
wire wadd1887d;
wire wadd1887c;
wire wadd1889d;
wire wadd1889c;
wire wadd1891d;
wire wadd1891c;
wire wadd1893d;
wire wadd1893c;
wire winv1895;
wire wboothprod1896;
wire wboothprod1897;
wire wboothprod1898;
wire wboothprod1899;
wire wcarry1900;
wire wcarry1901g;
wire wcarry1901p;
wire wcarry1903g;
wire wcarry1903p;
wire wcarry1905g;
wire wcarry1905p;
wire wcarry1907g;
wire wcarry1907p;
wire wadd1909d;
wire wadd1909c;
wire wadd1911d;
wire wadd1911c;
wire wadd1913d;
wire wadd1913c;
wire wadd1915d;
wire wadd1915c;
wire wboothprod1917;
wire wboothprod1918;
wire wboothprod1919;
wire wcarry1920;
wire wcarry1921g;
wire wcarry1921p;
wire wadd1923d;
wire wadd1923c;
wire wadd1925d;
wire wadd1925c;
wire wadd1927d;
wire wadd1927c;
wire winv1929;
wire wboothprod1930;
wire wboothprod1931;
wire wboothprod1932;
wire wcarry1933;
wire wcarry1934g;
wire wcarry1934p;
wire wcarry1936g;
wire wcarry1936p;
wire wadd1938d;
wire wadd1938c;
wire wadd1940d;
wire wadd1940c;
wire wadd1942d;
wire wadd1942c;
wire wboothprod1944;
wire wboothprod1945;
wire wcarry1946;
wire wcarry1947g;
wire wcarry1947p;
wire wadd1949d;
wire wadd1949c;
wire wadd1951d;
wire wadd1951c;
wire winv1953;
wire wboothprod1954;
wire wboothprod1955;
wire wcarry1956;
wire wcarry1957g;
wire wcarry1957p;
wire wcarry1959g;
wire wcarry1959p;
wire wcarry1961g;
wire wcarry1961p;
wire wadd1963d;
wire wadd1963c;
wire wadd1965d;
wire wadd1965c;
wire wboothprod1967;
wire wcarry1968;
wire wcarry1969g;
wire wcarry1969p;
wire wadd1971d;
wire wadd1971c;
wire winv1973;
wire wboothprod1974;
wire wcarry1975;
wire wcarry1976g;
wire wcarry1976p;
wire wcarry1978g;
wire wcarry1978p;
wire wadd1980d;
wire wadd1980c;
wire wcarry1982;
wire wcarry1983g;
wire wcarry1983p;
smul_booth_prod u0 ( 1'b0, x[0], x[1], 1'b0, y[0], wboothprod2 );
smul_booth_neg u1 ( 1'b0, x[0], x[1], wboothneg3 );
smul_full_add u2 ( wboothprod2, wboothneg3, 1'b0, wadd0d, wadd0c );
smul_booth_prod u3 ( 1'b0, x[0], x[1], y[0], y[1], wboothprod6 );
smul_carry_prop u4 ( wboothprod2, wboothneg3, wcarry8g, wcarry8p );
smul_carry_eval u5 ( wcarry8g, wcarry8p, 1'b0, wcarry7 );
smul_full_add u6 ( wboothprod6, 1'b0, wcarry7, wadd4d, wadd4c );
smul_booth_prod u7 ( 1'b0, x[0], x[1], y[1], y[2], wboothprod14 );
smul_booth_prod u8 ( x[1], x[2], x[3], 1'b0, y[0], wboothprod15 );
smul_booth_neg u9 ( x[1], x[2], x[3], wboothneg16 );
smul_full_add u10 ( wboothprod14, wboothprod15, wboothneg16, wadd12d, wadd12c );
smul_carry_prop u11 ( wboothprod6, 1'b0, wcarry20g, wcarry20p );
smul_carry_merge u12 ( wcarry8g, wcarry8p, wcarry20g, wcarry20p, wcarry18g, wcarry18p );
smul_carry_eval u13 ( wcarry18g, wcarry18p, 1'b0, wcarry17 );
smul_full_add u14 ( wadd12d, 1'b0, wcarry17, wadd10d, wadd10c );
smul_booth_prod u15 ( 1'b0, x[0], x[1], y[2], y[3], wboothprod26 );
smul_booth_prod u16 ( x[1], x[2], x[3], y[0], y[1], wboothprod27 );
smul_full_add u17 ( wadd12c, wboothprod26, wboothprod27, wadd24d, wadd24c );
smul_carry_prop u18 ( wadd12d, 1'b0, wcarry29g, wcarry29p );
smul_carry_eval u19 ( wcarry29g, wcarry29p, wcarry17, wcarry28 );
smul_full_add u20 ( wadd24d, 1'b0, wcarry28, wadd22d, wadd22c );
smul_booth_prod u21 ( 1'b0, x[0], x[1], y[3], y[4], wboothprod37 );
smul_booth_prod u22 ( x[1], x[2], x[3], y[1], y[2], wboothprod38 );
smul_booth_prod u23 ( x[3], x[4], x[5], 1'b0, y[0], wboothprod39 );
smul_full_add u24 ( wboothprod37, wboothprod38, wboothprod39, wadd35d, wadd35c );
smul_booth_neg u25 ( x[3], x[4], x[5], wboothneg40 );
smul_full_add u26 ( wadd24c, wadd35d, wboothneg40, wadd33d, wadd33c );
smul_carry_prop u27 ( wadd24d, 1'b0, wcarry46g, wcarry46p );
smul_carry_merge u28 ( wcarry29g, wcarry29p, wcarry46g, wcarry46p, wcarry44g, wcarry44p );
smul_carry_merge u29 ( wcarry18g, wcarry18p, wcarry44g, wcarry44p, wcarry42g, wcarry42p );
smul_carry_eval u30 ( wcarry42g, wcarry42p, 1'b0, wcarry41 );
smul_full_add u31 ( wadd33d, 1'b0, wcarry41, wadd31d, wadd31c );
smul_booth_prod u32 ( 1'b0, x[0], x[1], y[4], y[5], wboothprod54 );
smul_booth_prod u33 ( x[1], x[2], x[3], y[2], y[3], wboothprod55 );
smul_booth_prod u34 ( x[3], x[4], x[5], y[0], y[1], wboothprod56 );
smul_full_add u35 ( wboothprod54, wboothprod55, wboothprod56, wadd52d, wadd52c );
smul_full_add u36 ( wadd33c, wadd35c, wadd52d, wadd50d, wadd50c );
smul_carry_prop u37 ( wadd33d, 1'b0, wcarry58g, wcarry58p );
smul_carry_eval u38 ( wcarry58g, wcarry58p, wcarry41, wcarry57 );
smul_full_add u39 ( wadd50d, 1'b0, wcarry57, wadd48d, wadd48c );
smul_booth_prod u40 ( 1'b0, x[0], x[1], y[5], y[6], wboothprod66 );
smul_booth_prod u41 ( x[1], x[2], x[3], y[3], y[4], wboothprod67 );
smul_booth_prod u42 ( x[3], x[4], x[5], y[1], y[2], wboothprod68 );
smul_full_add u43 ( wboothprod66, wboothprod67, wboothprod68, wadd64d, wadd64c );
smul_booth_prod u44 ( x[5], x[6], x[7], 1'b0, y[0], wboothprod71 );
smul_booth_neg u45 ( x[5], x[6], x[7], wboothneg72 );
smul_half_add u46 ( wboothprod71, wboothneg72, wadd69d, wadd69c );
smul_full_add u47 ( wadd52c, wadd64d, wadd69d, wadd62d, wadd62c );
smul_carry_prop u48 ( wadd50d, 1'b0, wcarry76g, wcarry76p );
smul_carry_merge u49 ( wcarry58g, wcarry58p, wcarry76g, wcarry76p, wcarry74g, wcarry74p );
smul_carry_eval u50 ( wcarry74g, wcarry74p, wcarry41, wcarry73 );
smul_full_add u51 ( wadd50c, wadd62d, wcarry73, wadd60d, wadd60c );
smul_booth_prod u52 ( 1'b0, x[0], x[1], y[6], y[7], wboothprod86 );
smul_booth_prod u53 ( x[1], x[2], x[3], y[4], y[5], wboothprod87 );
smul_booth_prod u54 ( x[3], x[4], x[5], y[2], y[3], wboothprod88 );
smul_full_add u55 ( wboothprod86, wboothprod87, wboothprod88, wadd84d, wadd84c );
smul_full_add u56 ( wadd64c, wadd69c, wadd84d, wadd82d, wadd82c );
smul_booth_prod u57 ( x[5], x[6], x[7], y[0], y[1], wboothprod89 );
smul_full_add u58 ( wadd62c, wadd82d, wboothprod89, wadd80d, wadd80c );
smul_carry_prop u59 ( wadd50c, wadd62d, wcarry91g, wcarry91p );
smul_carry_eval u60 ( wcarry91g, wcarry91p, wcarry73, wcarry90 );
smul_full_add u61 ( wadd80d, 1'b0, wcarry90, wadd78d, wadd78c );
smul_booth_prod u62 ( 1'b0, x[0], x[1], y[7], y[8], wboothprod101 );
smul_booth_prod u63 ( x[1], x[2], x[3], y[5], y[6], wboothprod102 );
smul_booth_prod u64 ( x[3], x[4], x[5], y[3], y[4], wboothprod103 );
smul_full_add u65 ( wboothprod101, wboothprod102, wboothprod103, wadd99d, wadd99c );
smul_booth_prod u66 ( x[5], x[6], x[7], y[1], y[2], wboothprod106 );
smul_booth_prod u67 ( x[7], x[8], x[9], 1'b0, y[0], wboothprod107 );
smul_booth_neg u68 ( x[7], x[8], x[9], wboothneg108 );
smul_full_add u69 ( wboothprod106, wboothprod107, wboothneg108, wadd104d, wadd104c );
smul_full_add u70 ( wadd84c, wadd99d, wadd104d, wadd97d, wadd97c );
smul_full_add u71 ( wadd80c, wadd82c, wadd97d, wadd95d, wadd95c );
smul_carry_prop u72 ( wadd80d, 1'b0, wcarry116g, wcarry116p );
smul_carry_merge u73 ( wcarry91g, wcarry91p, wcarry116g, wcarry116p, wcarry114g, wcarry114p );
smul_carry_merge u74 ( wcarry74g, wcarry74p, wcarry114g, wcarry114p, wcarry112g, wcarry112p );
smul_carry_merge u75 ( wcarry42g, wcarry42p, wcarry112g, wcarry112p, wcarry110g, wcarry110p );
smul_carry_eval u76 ( wcarry110g, wcarry110p, 1'b0, wcarry109 );
smul_full_add u77 ( wadd95d, 1'b0, wcarry109, wadd93d, wadd93c );
smul_booth_prod u78 ( 1'b0, x[0], x[1], y[8], y[9], wboothprod126 );
smul_booth_prod u79 ( x[1], x[2], x[3], y[6], y[7], wboothprod127 );
smul_booth_prod u80 ( x[3], x[4], x[5], y[4], y[5], wboothprod128 );
smul_full_add u81 ( wboothprod126, wboothprod127, wboothprod128, wadd124d, wadd124c );
smul_full_add u82 ( wadd99c, wadd104c, wadd124d, wadd122d, wadd122c );
smul_booth_prod u83 ( x[5], x[6], x[7], y[2], y[3], wboothprod131 );
smul_booth_prod u84 ( x[7], x[8], x[9], y[0], y[1], wboothprod132 );
smul_half_add u85 ( wboothprod131, wboothprod132, wadd129d, wadd129c );
smul_full_add u86 ( wadd97c, wadd122d, wadd129d, wadd120d, wadd120c );
smul_carry_prop u87 ( wadd95d, 1'b0, wcarry134g, wcarry134p );
smul_carry_eval u88 ( wcarry134g, wcarry134p, wcarry109, wcarry133 );
smul_full_add u89 ( wadd95c, wadd120d, wcarry133, wadd118d, wadd118c );
smul_booth_prod u90 ( 1'b0, x[0], x[1], y[9], y[10], wboothprod146 );
smul_booth_prod u91 ( x[1], x[2], x[3], y[7], y[8], wboothprod147 );
smul_booth_prod u92 ( x[3], x[4], x[5], y[5], y[6], wboothprod148 );
smul_full_add u93 ( wboothprod146, wboothprod147, wboothprod148, wadd144d, wadd144c );
smul_booth_prod u94 ( x[5], x[6], x[7], y[3], y[4], wboothprod151 );
smul_booth_prod u95 ( x[7], x[8], x[9], y[1], y[2], wboothprod152 );
smul_booth_prod u96 ( x[9], x[10], x[11], 1'b0, y[0], wboothprod153 );
smul_full_add u97 ( wboothprod151, wboothprod152, wboothprod153, wadd149d, wadd149c );
smul_full_add u98 ( wadd124c, wadd144d, wadd149d, wadd142d, wadd142c );
smul_full_add u99 ( wadd122c, wadd129c, wadd142d, wadd140d, wadd140c );
smul_booth_neg u100 ( x[9], x[10], x[11], wboothneg154 );
smul_full_add u101 ( wadd120c, wadd140d, wboothneg154, wadd138d, wadd138c );
smul_carry_prop u102 ( wadd95c, wadd120d, wcarry158g, wcarry158p );
smul_carry_merge u103 ( wcarry134g, wcarry134p, wcarry158g, wcarry158p, wcarry156g, wcarry156p );
smul_carry_eval u104 ( wcarry156g, wcarry156p, wcarry109, wcarry155 );
smul_full_add u105 ( wadd138d, 1'b0, wcarry155, wadd136d, wadd136c );
smul_booth_prod u106 ( 1'b0, x[0], x[1], y[10], y[11], wboothprod170 );
smul_booth_prod u107 ( x[1], x[2], x[3], y[8], y[9], wboothprod171 );
smul_booth_prod u108 ( x[3], x[4], x[5], y[6], y[7], wboothprod172 );
smul_full_add u109 ( wboothprod170, wboothprod171, wboothprod172, wadd168d, wadd168c );
smul_full_add u110 ( wadd144c, wadd149c, wadd168d, wadd166d, wadd166c );
smul_booth_prod u111 ( x[5], x[6], x[7], y[4], y[5], wboothprod175 );
smul_booth_prod u112 ( x[7], x[8], x[9], y[2], y[3], wboothprod176 );
smul_booth_prod u113 ( x[9], x[10], x[11], y[0], y[1], wboothprod177 );
smul_full_add u114 ( wboothprod175, wboothprod176, wboothprod177, wadd173d, wadd173c );
smul_full_add u115 ( wadd142c, wadd166d, wadd173d, wadd164d, wadd164c );
smul_full_add u116 ( wadd138c, wadd140c, wadd164d, wadd162d, wadd162c );
smul_carry_prop u117 ( wadd138d, 1'b0, wcarry179g, wcarry179p );
smul_carry_eval u118 ( wcarry179g, wcarry179p, wcarry155, wcarry178 );
smul_full_add u119 ( wadd162d, 1'b0, wcarry178, wadd160d, wadd160c );
smul_booth_prod u120 ( 1'b0, x[0], x[1], y[11], y[12], wboothprod191 );
smul_booth_prod u121 ( x[1], x[2], x[3], y[9], y[10], wboothprod192 );
smul_booth_prod u122 ( x[3], x[4], x[5], y[7], y[8], wboothprod193 );
smul_full_add u123 ( wboothprod191, wboothprod192, wboothprod193, wadd189d, wadd189c );
smul_full_add u124 ( wadd168c, wadd173c, wadd189d, wadd187d, wadd187c );
smul_booth_prod u125 ( x[5], x[6], x[7], y[5], y[6], wboothprod198 );
smul_booth_prod u126 ( x[7], x[8], x[9], y[3], y[4], wboothprod199 );
smul_booth_prod u127 ( x[9], x[10], x[11], y[1], y[2], wboothprod200 );
smul_full_add u128 ( wboothprod198, wboothprod199, wboothprod200, wadd196d, wadd196c );
smul_booth_prod u129 ( x[11], x[12], x[13], 1'b0, y[0], wboothprod201 );
smul_booth_neg u130 ( x[11], x[12], x[13], wboothneg202 );
smul_full_add u131 ( wadd196d, wboothprod201, wboothneg202, wadd194d, wadd194c );
smul_full_add u132 ( wadd166c, wadd187d, wadd194d, wadd185d, wadd185c );
smul_full_add u133 ( wadd162c, wadd164c, wadd185d, wadd183d, wadd183c );
smul_carry_prop u134 ( wadd162d, 1'b0, wcarry208g, wcarry208p );
smul_carry_merge u135 ( wcarry179g, wcarry179p, wcarry208g, wcarry208p, wcarry206g, wcarry206p );
smul_carry_merge u136 ( wcarry156g, wcarry156p, wcarry206g, wcarry206p, wcarry204g, wcarry204p );
smul_carry_eval u137 ( wcarry204g, wcarry204p, wcarry109, wcarry203 );
smul_full_add u138 ( wadd183d, 1'b0, wcarry203, wadd181d, wadd181c );
smul_booth_prod u139 ( 1'b0, x[0], x[1], y[12], y[13], wboothprod220 );
smul_booth_prod u140 ( x[1], x[2], x[3], y[10], y[11], wboothprod221 );
smul_booth_prod u141 ( x[3], x[4], x[5], y[8], y[9], wboothprod222 );
smul_full_add u142 ( wboothprod220, wboothprod221, wboothprod222, wadd218d, wadd218c );
smul_full_add u143 ( wadd189c, wadd196c, wadd218d, wadd216d, wadd216c );
smul_full_add u144 ( wadd187c, wadd194c, wadd216d, wadd214d, wadd214c );
smul_booth_prod u145 ( x[5], x[6], x[7], y[6], y[7], wboothprod227 );
smul_booth_prod u146 ( x[7], x[8], x[9], y[4], y[5], wboothprod228 );
smul_booth_prod u147 ( x[9], x[10], x[11], y[2], y[3], wboothprod229 );
smul_full_add u148 ( wboothprod227, wboothprod228, wboothprod229, wadd225d, wadd225c );
smul_booth_prod u149 ( x[11], x[12], x[13], y[0], y[1], wboothprod230 );
smul_half_add u150 ( wadd225d, wboothprod230, wadd223d, wadd223c );
smul_full_add u151 ( wadd185c, wadd214d, wadd223d, wadd212d, wadd212c );
smul_carry_prop u152 ( wadd183d, 1'b0, wcarry232g, wcarry232p );
smul_carry_eval u153 ( wcarry232g, wcarry232p, wcarry203, wcarry231 );
smul_full_add u154 ( wadd183c, wadd212d, wcarry231, wadd210d, wadd210c );
smul_booth_prod u155 ( 1'b0, x[0], x[1], y[13], y[14], wboothprod244 );
smul_booth_prod u156 ( x[1], x[2], x[3], y[11], y[12], wboothprod245 );
smul_booth_prod u157 ( x[3], x[4], x[5], y[9], y[10], wboothprod246 );
smul_full_add u158 ( wboothprod244, wboothprod245, wboothprod246, wadd242d, wadd242c );
smul_full_add u159 ( wadd218c, wadd225c, wadd242d, wadd240d, wadd240c );
smul_booth_prod u160 ( x[5], x[6], x[7], y[7], y[8], wboothprod251 );
smul_booth_prod u161 ( x[7], x[8], x[9], y[5], y[6], wboothprod252 );
smul_booth_prod u162 ( x[9], x[10], x[11], y[3], y[4], wboothprod253 );
smul_full_add u163 ( wboothprod251, wboothprod252, wboothprod253, wadd249d, wadd249c );
smul_booth_prod u164 ( x[11], x[12], x[13], y[1], y[2], wboothprod256 );
smul_booth_prod u165 ( x[13], x[14], x[15], 1'b0, y[0], wboothprod257 );
smul_booth_neg u166 ( x[13], x[14], x[15], wboothneg258 );
smul_full_add u167 ( wboothprod256, wboothprod257, wboothneg258, wadd254d, wadd254c );
smul_half_add u168 ( wadd249d, wadd254d, wadd247d, wadd247c );
smul_full_add u169 ( wadd216c, wadd240d, wadd247d, wadd238d, wadd238c );
smul_full_add u170 ( wadd214c, wadd223c, wadd238d, wadd236d, wadd236c );
smul_carry_prop u171 ( wadd183c, wadd212d, wcarry262g, wcarry262p );
smul_carry_merge u172 ( wcarry232g, wcarry232p, wcarry262g, wcarry262p, wcarry260g, wcarry260p );
smul_carry_eval u173 ( wcarry260g, wcarry260p, wcarry203, wcarry259 );
smul_full_add u174 ( wadd212c, wadd236d, wcarry259, wadd234d, wadd234c );
smul_full_add u175 ( wadd242c, wadd249c, wadd254c, wadd270d, wadd270c );
smul_full_add u176 ( wadd240c, wadd247c, wadd270d, wadd268d, wadd268c );
smul_booth_prod u177 ( 1'b0, x[0], x[1], y[14], y[15], wboothprod276 );
smul_booth_prod u178 ( x[1], x[2], x[3], y[12], y[13], wboothprod277 );
smul_booth_prod u179 ( x[3], x[4], x[5], y[10], y[11], wboothprod278 );
smul_full_add u180 ( wboothprod276, wboothprod277, wboothprod278, wadd274d, wadd274c );
smul_booth_prod u181 ( x[5], x[6], x[7], y[8], y[9], wboothprod281 );
smul_booth_prod u182 ( x[7], x[8], x[9], y[6], y[7], wboothprod282 );
smul_booth_prod u183 ( x[9], x[10], x[11], y[4], y[5], wboothprod283 );
smul_full_add u184 ( wboothprod281, wboothprod282, wboothprod283, wadd279d, wadd279c );
smul_booth_prod u185 ( x[11], x[12], x[13], y[2], y[3], wboothprod286 );
smul_booth_prod u186 ( x[13], x[14], x[15], y[0], y[1], wboothprod287 );
smul_half_add u187 ( wboothprod286, wboothprod287, wadd284d, wadd284c );
smul_full_add u188 ( wadd274d, wadd279d, wadd284d, wadd272d, wadd272c );
smul_full_add u189 ( wadd238c, wadd268d, wadd272d, wadd266d, wadd266c );
smul_carry_prop u190 ( wadd212c, wadd236d, wcarry289g, wcarry289p );
smul_carry_eval u191 ( wcarry289g, wcarry289p, wcarry259, wcarry288 );
smul_full_add u192 ( wadd236c, wadd266d, wcarry288, wadd264d, wadd264c );
smul_full_add u193 ( wadd274c, wadd279c, wadd284c, wadd297d, wadd297c );
smul_full_add u194 ( wadd270c, wadd272c, wadd297d, wadd295d, wadd295c );
smul_booth_prod u195 ( 1'b0, x[0], x[1], y[15], y[16], wboothprod305 );
smul_booth_prod u196 ( x[1], x[2], x[3], y[13], y[14], wboothprod306 );
smul_booth_prod u197 ( x[3], x[4], x[5], y[11], y[12], wboothprod307 );
smul_full_add u198 ( wboothprod305, wboothprod306, wboothprod307, wadd303d, wadd303c );
smul_booth_prod u199 ( x[5], x[6], x[7], y[9], y[10], wboothprod310 );
smul_booth_prod u200 ( x[7], x[8], x[9], y[7], y[8], wboothprod311 );
smul_booth_prod u201 ( x[9], x[10], x[11], y[5], y[6], wboothprod312 );
smul_full_add u202 ( wboothprod310, wboothprod311, wboothprod312, wadd308d, wadd308c );
smul_booth_prod u203 ( x[11], x[12], x[13], y[3], y[4], wboothprod315 );
smul_booth_prod u204 ( x[13], x[14], x[15], y[1], y[2], wboothprod316 );
smul_booth_prod u205 ( x[15], x[16], x[17], 1'b0, y[0], wboothprod317 );
smul_full_add u206 ( wboothprod315, wboothprod316, wboothprod317, wadd313d, wadd313c );
smul_full_add u207 ( wadd303d, wadd308d, wadd313d, wadd301d, wadd301c );
smul_booth_neg u208 ( x[15], x[16], x[17], wboothneg318 );
smul_half_add u209 ( wadd301d, wboothneg318, wadd299d, wadd299c );
smul_full_add u210 ( wadd268c, wadd295d, wadd299d, wadd293d, wadd293c );
smul_carry_prop u211 ( wadd236c, wadd266d, wcarry328g, wcarry328p );
smul_carry_merge u212 ( wcarry289g, wcarry289p, wcarry328g, wcarry328p, wcarry326g, wcarry326p );
smul_carry_merge u213 ( wcarry260g, wcarry260p, wcarry326g, wcarry326p, wcarry324g, wcarry324p );
smul_carry_merge u214 ( wcarry204g, wcarry204p, wcarry324g, wcarry324p, wcarry322g, wcarry322p );
smul_carry_merge u215 ( wcarry110g, wcarry110p, wcarry322g, wcarry322p, wcarry320g, wcarry320p );
smul_carry_eval u216 ( wcarry320g, wcarry320p, 1'b0, wcarry319 );
smul_full_add u217 ( wadd266c, wadd293d, wcarry319, wadd291d, wadd291c );
smul_full_add u218 ( wadd303c, wadd308c, wadd313c, wadd338d, wadd338c );
smul_full_add u219 ( wadd297c, wadd301c, wadd338d, wadd336d, wadd336c );
smul_full_add u220 ( wadd295c, wadd299c, wadd336d, wadd334d, wadd334c );
smul_booth_prod u221 ( 1'b0, x[0], x[1], y[16], y[17], wboothprod344 );
smul_booth_prod u222 ( x[1], x[2], x[3], y[14], y[15], wboothprod345 );
smul_booth_prod u223 ( x[3], x[4], x[5], y[12], y[13], wboothprod346 );
smul_full_add u224 ( wboothprod344, wboothprod345, wboothprod346, wadd342d, wadd342c );
smul_booth_prod u225 ( x[5], x[6], x[7], y[10], y[11], wboothprod349 );
smul_booth_prod u226 ( x[7], x[8], x[9], y[8], y[9], wboothprod350 );
smul_booth_prod u227 ( x[9], x[10], x[11], y[6], y[7], wboothprod351 );
smul_full_add u228 ( wboothprod349, wboothprod350, wboothprod351, wadd347d, wadd347c );
smul_booth_prod u229 ( x[11], x[12], x[13], y[4], y[5], wboothprod354 );
smul_booth_prod u230 ( x[13], x[14], x[15], y[2], y[3], wboothprod355 );
smul_booth_prod u231 ( x[15], x[16], x[17], y[0], y[1], wboothprod356 );
smul_full_add u232 ( wboothprod354, wboothprod355, wboothprod356, wadd352d, wadd352c );
smul_full_add u233 ( wadd342d, wadd347d, wadd352d, wadd340d, wadd340c );
smul_full_add u234 ( wadd293c, wadd334d, wadd340d, wadd332d, wadd332c );
smul_carry_prop u235 ( wadd266c, wadd293d, wcarry358g, wcarry358p );
smul_carry_eval u236 ( wcarry358g, wcarry358p, wcarry319, wcarry357 );
smul_full_add u237 ( wadd332d, 1'b0, wcarry357, wadd330d, wadd330c );
smul_full_add u238 ( wadd342c, wadd347c, wadd352c, wadd368d, wadd368c );
smul_full_add u239 ( wadd338c, wadd340c, wadd368d, wadd366d, wadd366c );
smul_booth_prod u240 ( 1'b0, x[0], x[1], y[17], y[18], wboothprod376 );
smul_booth_prod u241 ( x[1], x[2], x[3], y[15], y[16], wboothprod377 );
smul_booth_prod u242 ( x[3], x[4], x[5], y[13], y[14], wboothprod378 );
smul_full_add u243 ( wboothprod376, wboothprod377, wboothprod378, wadd374d, wadd374c );
smul_booth_prod u244 ( x[5], x[6], x[7], y[11], y[12], wboothprod381 );
smul_booth_prod u245 ( x[7], x[8], x[9], y[9], y[10], wboothprod382 );
smul_booth_prod u246 ( x[9], x[10], x[11], y[7], y[8], wboothprod383 );
smul_full_add u247 ( wboothprod381, wboothprod382, wboothprod383, wadd379d, wadd379c );
smul_booth_prod u248 ( x[11], x[12], x[13], y[5], y[6], wboothprod386 );
smul_booth_prod u249 ( x[13], x[14], x[15], y[3], y[4], wboothprod387 );
smul_booth_prod u250 ( x[15], x[16], x[17], y[1], y[2], wboothprod388 );
smul_full_add u251 ( wboothprod386, wboothprod387, wboothprod388, wadd384d, wadd384c );
smul_full_add u252 ( wadd374d, wadd379d, wadd384d, wadd372d, wadd372c );
smul_booth_prod u253 ( x[17], x[18], x[19], 1'b0, y[0], wboothprod389 );
smul_booth_neg u254 ( x[17], x[18], x[19], wboothneg390 );
smul_full_add u255 ( wadd372d, wboothprod389, wboothneg390, wadd370d, wadd370c );
smul_full_add u256 ( wadd336c, wadd366d, wadd370d, wadd364d, wadd364c );
smul_full_add u257 ( wadd332c, wadd334c, wadd364d, wadd362d, wadd362c );
smul_carry_prop u258 ( wadd332d, 1'b0, wcarry394g, wcarry394p );
smul_carry_merge u259 ( wcarry358g, wcarry358p, wcarry394g, wcarry394p, wcarry392g, wcarry392p );
smul_carry_eval u260 ( wcarry392g, wcarry392p, wcarry319, wcarry391 );
smul_full_add u261 ( wadd362d, 1'b0, wcarry391, wadd360d, wadd360c );
smul_full_add u262 ( wadd374c, wadd379c, wadd384c, wadd404d, wadd404c );
smul_full_add u263 ( wadd368c, wadd372c, wadd404d, wadd402d, wadd402c );
smul_full_add u264 ( wadd366c, wadd370c, wadd402d, wadd400d, wadd400c );
smul_booth_prod u265 ( 1'b0, x[0], x[1], y[18], y[19], wboothprod412 );
smul_booth_prod u266 ( x[1], x[2], x[3], y[16], y[17], wboothprod413 );
smul_booth_prod u267 ( x[3], x[4], x[5], y[14], y[15], wboothprod414 );
smul_full_add u268 ( wboothprod412, wboothprod413, wboothprod414, wadd410d, wadd410c );
smul_booth_prod u269 ( x[5], x[6], x[7], y[12], y[13], wboothprod417 );
smul_booth_prod u270 ( x[7], x[8], x[9], y[10], y[11], wboothprod418 );
smul_booth_prod u271 ( x[9], x[10], x[11], y[8], y[9], wboothprod419 );
smul_full_add u272 ( wboothprod417, wboothprod418, wboothprod419, wadd415d, wadd415c );
smul_booth_prod u273 ( x[11], x[12], x[13], y[6], y[7], wboothprod422 );
smul_booth_prod u274 ( x[13], x[14], x[15], y[4], y[5], wboothprod423 );
smul_booth_prod u275 ( x[15], x[16], x[17], y[2], y[3], wboothprod424 );
smul_full_add u276 ( wboothprod422, wboothprod423, wboothprod424, wadd420d, wadd420c );
smul_full_add u277 ( wadd410d, wadd415d, wadd420d, wadd408d, wadd408c );
smul_booth_prod u278 ( x[17], x[18], x[19], y[0], y[1], wboothprod425 );
smul_half_add u279 ( wadd408d, wboothprod425, wadd406d, wadd406c );
smul_full_add u280 ( wadd364c, wadd400d, wadd406d, wadd398d, wadd398c );
smul_carry_prop u281 ( wadd362d, 1'b0, wcarry427g, wcarry427p );
smul_carry_eval u282 ( wcarry427g, wcarry427p, wcarry391, wcarry426 );
smul_full_add u283 ( wadd362c, wadd398d, wcarry426, wadd396d, wadd396c );
smul_full_add u284 ( wadd410c, wadd415c, wadd420c, wadd437d, wadd437c );
smul_full_add u285 ( wadd404c, wadd408c, wadd437d, wadd435d, wadd435c );
smul_booth_prod u286 ( 1'b0, x[0], x[1], y[19], y[20], wboothprod445 );
smul_booth_prod u287 ( x[1], x[2], x[3], y[17], y[18], wboothprod446 );
smul_booth_prod u288 ( x[3], x[4], x[5], y[15], y[16], wboothprod447 );
smul_full_add u289 ( wboothprod445, wboothprod446, wboothprod447, wadd443d, wadd443c );
smul_booth_prod u290 ( x[5], x[6], x[7], y[13], y[14], wboothprod450 );
smul_booth_prod u291 ( x[7], x[8], x[9], y[11], y[12], wboothprod451 );
smul_booth_prod u292 ( x[9], x[10], x[11], y[9], y[10], wboothprod452 );
smul_full_add u293 ( wboothprod450, wboothprod451, wboothprod452, wadd448d, wadd448c );
smul_booth_prod u294 ( x[11], x[12], x[13], y[7], y[8], wboothprod455 );
smul_booth_prod u295 ( x[13], x[14], x[15], y[5], y[6], wboothprod456 );
smul_booth_prod u296 ( x[15], x[16], x[17], y[3], y[4], wboothprod457 );
smul_full_add u297 ( wboothprod455, wboothprod456, wboothprod457, wadd453d, wadd453c );
smul_full_add u298 ( wadd443d, wadd448d, wadd453d, wadd441d, wadd441c );
smul_booth_prod u299 ( x[17], x[18], x[19], y[1], y[2], wboothprod460 );
smul_booth_prod u300 ( x[19], x[20], x[21], 1'b0, y[0], wboothprod461 );
smul_booth_neg u301 ( x[19], x[20], x[21], wboothneg462 );
smul_full_add u302 ( wboothprod460, wboothprod461, wboothneg462, wadd458d, wadd458c );
smul_half_add u303 ( wadd441d, wadd458d, wadd439d, wadd439c );
smul_full_add u304 ( wadd402c, wadd435d, wadd439d, wadd433d, wadd433c );
smul_full_add u305 ( wadd400c, wadd406c, wadd433d, wadd431d, wadd431c );
smul_carry_prop u306 ( wadd362c, wadd398d, wcarry468g, wcarry468p );
smul_carry_merge u307 ( wcarry427g, wcarry427p, wcarry468g, wcarry468p, wcarry466g, wcarry466p );
smul_carry_merge u308 ( wcarry392g, wcarry392p, wcarry466g, wcarry466p, wcarry464g, wcarry464p );
smul_carry_eval u309 ( wcarry464g, wcarry464p, wcarry319, wcarry463 );
smul_full_add u310 ( wadd398c, wadd431d, wcarry463, wadd429d, wadd429c );
smul_full_add u311 ( wadd443c, wadd448c, wadd453c, wadd478d, wadd478c );
smul_full_add u312 ( wadd437c, wadd441c, wadd478d, wadd476d, wadd476c );
smul_full_add u313 ( wadd435c, wadd439c, wadd476d, wadd474d, wadd474c );
smul_booth_prod u314 ( 1'b0, x[0], x[1], y[20], y[21], wboothprod486 );
smul_booth_prod u315 ( x[1], x[2], x[3], y[18], y[19], wboothprod487 );
smul_booth_prod u316 ( x[3], x[4], x[5], y[16], y[17], wboothprod488 );
smul_full_add u317 ( wboothprod486, wboothprod487, wboothprod488, wadd484d, wadd484c );
smul_booth_prod u318 ( x[5], x[6], x[7], y[14], y[15], wboothprod491 );
smul_booth_prod u319 ( x[7], x[8], x[9], y[12], y[13], wboothprod492 );
smul_booth_prod u320 ( x[9], x[10], x[11], y[10], y[11], wboothprod493 );
smul_full_add u321 ( wboothprod491, wboothprod492, wboothprod493, wadd489d, wadd489c );
smul_full_add u322 ( wadd458c, wadd484d, wadd489d, wadd482d, wadd482c );
smul_booth_prod u323 ( x[11], x[12], x[13], y[8], y[9], wboothprod498 );
smul_booth_prod u324 ( x[13], x[14], x[15], y[6], y[7], wboothprod499 );
smul_booth_prod u325 ( x[15], x[16], x[17], y[4], y[5], wboothprod500 );
smul_full_add u326 ( wboothprod498, wboothprod499, wboothprod500, wadd496d, wadd496c );
smul_booth_prod u327 ( x[17], x[18], x[19], y[2], y[3], wboothprod501 );
smul_booth_prod u328 ( x[19], x[20], x[21], y[0], y[1], wboothprod502 );
smul_full_add u329 ( wadd496d, wboothprod501, wboothprod502, wadd494d, wadd494c );
smul_half_add u330 ( wadd482d, wadd494d, wadd480d, wadd480c );
smul_full_add u331 ( wadd433c, wadd474d, wadd480d, wadd472d, wadd472c );
smul_carry_prop u332 ( wadd398c, wadd431d, wcarry504g, wcarry504p );
smul_carry_eval u333 ( wcarry504g, wcarry504p, wcarry463, wcarry503 );
smul_full_add u334 ( wadd431c, wadd472d, wcarry503, wadd470d, wadd470c );
smul_full_add u335 ( wadd478c, wadd482c, wadd494c, wadd512d, wadd512c );
smul_full_add u336 ( wadd484c, wadd489c, wadd496c, wadd516d, wadd516c );
smul_booth_prod u337 ( 1'b0, x[0], x[1], y[21], y[22], wboothprod522 );
smul_booth_prod u338 ( x[1], x[2], x[3], y[19], y[20], wboothprod523 );
smul_booth_prod u339 ( x[3], x[4], x[5], y[17], y[18], wboothprod524 );
smul_full_add u340 ( wboothprod522, wboothprod523, wboothprod524, wadd520d, wadd520c );
smul_booth_prod u341 ( x[5], x[6], x[7], y[15], y[16], wboothprod527 );
smul_booth_prod u342 ( x[7], x[8], x[9], y[13], y[14], wboothprod528 );
smul_booth_prod u343 ( x[9], x[10], x[11], y[11], y[12], wboothprod529 );
smul_full_add u344 ( wboothprod527, wboothprod528, wboothprod529, wadd525d, wadd525c );
smul_booth_prod u345 ( x[11], x[12], x[13], y[9], y[10], wboothprod532 );
smul_booth_prod u346 ( x[13], x[14], x[15], y[7], y[8], wboothprod533 );
smul_booth_prod u347 ( x[15], x[16], x[17], y[5], y[6], wboothprod534 );
smul_full_add u348 ( wboothprod532, wboothprod533, wboothprod534, wadd530d, wadd530c );
smul_full_add u349 ( wadd520d, wadd525d, wadd530d, wadd518d, wadd518c );
smul_booth_prod u350 ( x[17], x[18], x[19], y[3], y[4], wboothprod539 );
smul_booth_prod u351 ( x[19], x[20], x[21], y[1], y[2], wboothprod540 );
smul_booth_prod u352 ( x[21], x[22], x[23], 1'b0, y[0], wboothprod541 );
smul_full_add u353 ( wboothprod539, wboothprod540, wboothprod541, wadd537d, wadd537c );
smul_booth_neg u354 ( x[21], x[22], x[23], wboothneg542 );
smul_half_add u355 ( wadd537d, wboothneg542, wadd535d, wadd535c );
smul_full_add u356 ( wadd516d, wadd518d, wadd535d, wadd514d, wadd514c );
smul_full_add u357 ( wadd476c, wadd512d, wadd514d, wadd510d, wadd510c );
smul_full_add u358 ( wadd474c, wadd480c, wadd510d, wadd508d, wadd508c );
smul_carry_prop u359 ( wadd431c, wadd472d, wcarry546g, wcarry546p );
smul_carry_merge u360 ( wcarry504g, wcarry504p, wcarry546g, wcarry546p, wcarry544g, wcarry544p );
smul_carry_eval u361 ( wcarry544g, wcarry544p, wcarry463, wcarry543 );
smul_full_add u362 ( wadd472c, wadd508d, wcarry543, wadd506d, wadd506c );
smul_full_add u363 ( wadd516c, wadd518c, wadd535c, wadd554d, wadd554c );
smul_full_add u364 ( wadd512c, wadd514c, wadd554d, wadd552d, wadd552c );
smul_full_add u365 ( wadd520c, wadd525c, wadd530c, wadd558d, wadd558c );
smul_booth_prod u366 ( 1'b0, x[0], x[1], y[22], y[23], wboothprod564 );
smul_booth_prod u367 ( x[1], x[2], x[3], y[20], y[21], wboothprod565 );
smul_booth_prod u368 ( x[3], x[4], x[5], y[18], y[19], wboothprod566 );
smul_full_add u369 ( wboothprod564, wboothprod565, wboothprod566, wadd562d, wadd562c );
smul_booth_prod u370 ( x[5], x[6], x[7], y[16], y[17], wboothprod569 );
smul_booth_prod u371 ( x[7], x[8], x[9], y[14], y[15], wboothprod570 );
smul_booth_prod u372 ( x[9], x[10], x[11], y[12], y[13], wboothprod571 );
smul_full_add u373 ( wboothprod569, wboothprod570, wboothprod571, wadd567d, wadd567c );
smul_full_add u374 ( wadd537c, wadd562d, wadd567d, wadd560d, wadd560c );
smul_booth_prod u375 ( x[11], x[12], x[13], y[10], y[11], wboothprod576 );
smul_booth_prod u376 ( x[13], x[14], x[15], y[8], y[9], wboothprod577 );
smul_booth_prod u377 ( x[15], x[16], x[17], y[6], y[7], wboothprod578 );
smul_full_add u378 ( wboothprod576, wboothprod577, wboothprod578, wadd574d, wadd574c );
smul_booth_prod u379 ( x[17], x[18], x[19], y[4], y[5], wboothprod581 );
smul_booth_prod u380 ( x[19], x[20], x[21], y[2], y[3], wboothprod582 );
smul_booth_prod u381 ( x[21], x[22], x[23], y[0], y[1], wboothprod583 );
smul_full_add u382 ( wboothprod581, wboothprod582, wboothprod583, wadd579d, wadd579c );
smul_half_add u383 ( wadd574d, wadd579d, wadd572d, wadd572c );
smul_full_add u384 ( wadd558d, wadd560d, wadd572d, wadd556d, wadd556c );
smul_full_add u385 ( wadd510c, wadd552d, wadd556d, wadd550d, wadd550c );
smul_carry_prop u386 ( wadd472c, wadd508d, wcarry585g, wcarry585p );
smul_carry_eval u387 ( wcarry585g, wcarry585p, wcarry543, wcarry584 );
smul_full_add u388 ( wadd508c, wadd550d, wcarry584, wadd548d, wadd548c );
smul_full_add u389 ( wadd558c, wadd560c, wadd572c, wadd593d, wadd593c );
smul_full_add u390 ( wadd554c, wadd556c, wadd593d, wadd591d, wadd591c );
smul_full_add u391 ( wadd562c, wadd567c, wadd574c, wadd597d, wadd597c );
smul_booth_prod u392 ( 1'b0, x[0], x[1], y[23], y[24], wboothprod603 );
smul_booth_prod u393 ( x[1], x[2], x[3], y[21], y[22], wboothprod604 );
smul_booth_prod u394 ( x[3], x[4], x[5], y[19], y[20], wboothprod605 );
smul_full_add u395 ( wboothprod603, wboothprod604, wboothprod605, wadd601d, wadd601c );
smul_booth_prod u396 ( x[5], x[6], x[7], y[17], y[18], wboothprod608 );
smul_booth_prod u397 ( x[7], x[8], x[9], y[15], y[16], wboothprod609 );
smul_booth_prod u398 ( x[9], x[10], x[11], y[13], y[14], wboothprod610 );
smul_full_add u399 ( wboothprod608, wboothprod609, wboothprod610, wadd606d, wadd606c );
smul_full_add u400 ( wadd579c, wadd601d, wadd606d, wadd599d, wadd599c );
smul_booth_prod u401 ( x[11], x[12], x[13], y[11], y[12], wboothprod615 );
smul_booth_prod u402 ( x[13], x[14], x[15], y[9], y[10], wboothprod616 );
smul_booth_prod u403 ( x[15], x[16], x[17], y[7], y[8], wboothprod617 );
smul_full_add u404 ( wboothprod615, wboothprod616, wboothprod617, wadd613d, wadd613c );
smul_booth_prod u405 ( x[17], x[18], x[19], y[5], y[6], wboothprod620 );
smul_booth_prod u406 ( x[19], x[20], x[21], y[3], y[4], wboothprod621 );
smul_booth_prod u407 ( x[21], x[22], x[23], y[1], y[2], wboothprod622 );
smul_full_add u408 ( wboothprod620, wboothprod621, wboothprod622, wadd618d, wadd618c );
smul_booth_prod u409 ( x[23], x[24], x[25], 1'b0, y[0], wboothprod625 );
smul_booth_neg u410 ( x[23], x[24], x[25], wboothneg626 );
smul_half_add u411 ( wboothprod625, wboothneg626, wadd623d, wadd623c );
smul_full_add u412 ( wadd613d, wadd618d, wadd623d, wadd611d, wadd611c );
smul_full_add u413 ( wadd597d, wadd599d, wadd611d, wadd595d, wadd595c );
smul_full_add u414 ( wadd552c, wadd591d, wadd595d, wadd589d, wadd589c );
smul_carry_prop u415 ( wadd508c, wadd550d, wcarry634g, wcarry634p );
smul_carry_merge u416 ( wcarry585g, wcarry585p, wcarry634g, wcarry634p, wcarry632g, wcarry632p );
smul_carry_merge u417 ( wcarry544g, wcarry544p, wcarry632g, wcarry632p, wcarry630g, wcarry630p );
smul_carry_merge u418 ( wcarry464g, wcarry464p, wcarry630g, wcarry630p, wcarry628g, wcarry628p );
smul_carry_eval u419 ( wcarry628g, wcarry628p, wcarry319, wcarry627 );
smul_full_add u420 ( wadd550c, wadd589d, wcarry627, wadd587d, wadd587c );
smul_full_add u421 ( wadd597c, wadd599c, wadd611c, wadd642d, wadd642c );
smul_full_add u422 ( wadd593c, wadd595c, wadd642d, wadd640d, wadd640c );
smul_full_add u423 ( wadd601c, wadd606c, wadd613c, wadd648d, wadd648c );
smul_booth_prod u424 ( 1'b0, x[0], x[1], y[24], y[25], wboothprod654 );
smul_booth_prod u425 ( x[1], x[2], x[3], y[22], y[23], wboothprod655 );
smul_booth_prod u426 ( x[3], x[4], x[5], y[20], y[21], wboothprod656 );
smul_full_add u427 ( wboothprod654, wboothprod655, wboothprod656, wadd652d, wadd652c );
smul_full_add u428 ( wadd618c, wadd623c, wadd652d, wadd650d, wadd650c );
smul_booth_prod u429 ( x[5], x[6], x[7], y[18], y[19], wboothprod661 );
smul_booth_prod u430 ( x[7], x[8], x[9], y[16], y[17], wboothprod662 );
smul_booth_prod u431 ( x[9], x[10], x[11], y[14], y[15], wboothprod663 );
smul_full_add u432 ( wboothprod661, wboothprod662, wboothprod663, wadd659d, wadd659c );
smul_booth_prod u433 ( x[11], x[12], x[13], y[12], y[13], wboothprod666 );
smul_booth_prod u434 ( x[13], x[14], x[15], y[10], y[11], wboothprod667 );
smul_booth_prod u435 ( x[15], x[16], x[17], y[8], y[9], wboothprod668 );
smul_full_add u436 ( wboothprod666, wboothprod667, wboothprod668, wadd664d, wadd664c );
smul_booth_prod u437 ( x[17], x[18], x[19], y[6], y[7], wboothprod671 );
smul_booth_prod u438 ( x[19], x[20], x[21], y[4], y[5], wboothprod672 );
smul_booth_prod u439 ( x[21], x[22], x[23], y[2], y[3], wboothprod673 );
smul_full_add u440 ( wboothprod671, wboothprod672, wboothprod673, wadd669d, wadd669c );
smul_full_add u441 ( wadd659d, wadd664d, wadd669d, wadd657d, wadd657c );
smul_full_add u442 ( wadd648d, wadd650d, wadd657d, wadd646d, wadd646c );
smul_booth_prod u443 ( x[23], x[24], x[25], y[0], y[1], wboothprod674 );
smul_half_add u444 ( wadd646d, wboothprod674, wadd644d, wadd644c );
smul_full_add u445 ( wadd591c, wadd640d, wadd644d, wadd638d, wadd638c );
smul_carry_prop u446 ( wadd550c, wadd589d, wcarry676g, wcarry676p );
smul_carry_eval u447 ( wcarry676g, wcarry676p, wcarry627, wcarry675 );
smul_full_add u448 ( wadd589c, wadd638d, wcarry675, wadd636d, wadd636c );
smul_full_add u449 ( wadd648c, wadd650c, wadd657c, wadd686d, wadd686c );
smul_full_add u450 ( wadd642c, wadd646c, wadd686d, wadd684d, wadd684c );
smul_full_add u451 ( wadd640c, wadd644c, wadd684d, wadd682d, wadd682c );
smul_full_add u452 ( wadd652c, wadd659c, wadd664c, wadd690d, wadd690c );
smul_booth_prod u453 ( 1'b0, x[0], x[1], y[25], y[26], wboothprod696 );
smul_booth_prod u454 ( x[1], x[2], x[3], y[23], y[24], wboothprod697 );
smul_booth_prod u455 ( x[3], x[4], x[5], y[21], y[22], wboothprod698 );
smul_full_add u456 ( wboothprod696, wboothprod697, wboothprod698, wadd694d, wadd694c );
smul_booth_prod u457 ( x[5], x[6], x[7], y[19], y[20], wboothprod701 );
smul_booth_prod u458 ( x[7], x[8], x[9], y[17], y[18], wboothprod702 );
smul_booth_prod u459 ( x[9], x[10], x[11], y[15], y[16], wboothprod703 );
smul_full_add u460 ( wboothprod701, wboothprod702, wboothprod703, wadd699d, wadd699c );
smul_full_add u461 ( wadd669c, wadd694d, wadd699d, wadd692d, wadd692c );
smul_booth_prod u462 ( x[11], x[12], x[13], y[13], y[14], wboothprod708 );
smul_booth_prod u463 ( x[13], x[14], x[15], y[11], y[12], wboothprod709 );
smul_booth_prod u464 ( x[15], x[16], x[17], y[9], y[10], wboothprod710 );
smul_full_add u465 ( wboothprod708, wboothprod709, wboothprod710, wadd706d, wadd706c );
smul_booth_prod u466 ( x[17], x[18], x[19], y[7], y[8], wboothprod713 );
smul_booth_prod u467 ( x[19], x[20], x[21], y[5], y[6], wboothprod714 );
smul_booth_prod u468 ( x[21], x[22], x[23], y[3], y[4], wboothprod715 );
smul_full_add u469 ( wboothprod713, wboothprod714, wboothprod715, wadd711d, wadd711c );
smul_booth_prod u470 ( x[23], x[24], x[25], y[1], y[2], wboothprod718 );
smul_booth_prod u471 ( x[25], x[26], x[27], 1'b0, y[0], wboothprod719 );
smul_booth_neg u472 ( x[25], x[26], x[27], wboothneg720 );
smul_full_add u473 ( wboothprod718, wboothprod719, wboothneg720, wadd716d, wadd716c );
smul_full_add u474 ( wadd706d, wadd711d, wadd716d, wadd704d, wadd704c );
smul_full_add u475 ( wadd690d, wadd692d, wadd704d, wadd688d, wadd688c );
smul_full_add u476 ( wadd638c, wadd682d, wadd688d, wadd680d, wadd680c );
smul_carry_prop u477 ( wadd589c, wadd638d, wcarry724g, wcarry724p );
smul_carry_merge u478 ( wcarry676g, wcarry676p, wcarry724g, wcarry724p, wcarry722g, wcarry722p );
smul_carry_eval u479 ( wcarry722g, wcarry722p, wcarry627, wcarry721 );
smul_full_add u480 ( wadd680d, 1'b0, wcarry721, wadd678d, wadd678c );
smul_full_add u481 ( wadd690c, wadd692c, wadd704c, wadd734d, wadd734c );
smul_full_add u482 ( wadd686c, wadd688c, wadd734d, wadd732d, wadd732c );
smul_full_add u483 ( wadd694c, wadd699c, wadd706c, wadd740d, wadd740c );
smul_booth_prod u484 ( 1'b0, x[0], x[1], y[26], y[27], wboothprod746 );
smul_booth_prod u485 ( x[1], x[2], x[3], y[24], y[25], wboothprod747 );
smul_booth_prod u486 ( x[3], x[4], x[5], y[22], y[23], wboothprod748 );
smul_full_add u487 ( wboothprod746, wboothprod747, wboothprod748, wadd744d, wadd744c );
smul_full_add u488 ( wadd711c, wadd716c, wadd744d, wadd742d, wadd742c );
smul_booth_prod u489 ( x[5], x[6], x[7], y[20], y[21], wboothprod753 );
smul_booth_prod u490 ( x[7], x[8], x[9], y[18], y[19], wboothprod754 );
smul_booth_prod u491 ( x[9], x[10], x[11], y[16], y[17], wboothprod755 );
smul_full_add u492 ( wboothprod753, wboothprod754, wboothprod755, wadd751d, wadd751c );
smul_booth_prod u493 ( x[11], x[12], x[13], y[14], y[15], wboothprod758 );
smul_booth_prod u494 ( x[13], x[14], x[15], y[12], y[13], wboothprod759 );
smul_booth_prod u495 ( x[15], x[16], x[17], y[10], y[11], wboothprod760 );
smul_full_add u496 ( wboothprod758, wboothprod759, wboothprod760, wadd756d, wadd756c );
smul_booth_prod u497 ( x[17], x[18], x[19], y[8], y[9], wboothprod763 );
smul_booth_prod u498 ( x[19], x[20], x[21], y[6], y[7], wboothprod764 );
smul_booth_prod u499 ( x[21], x[22], x[23], y[4], y[5], wboothprod765 );
smul_full_add u500 ( wboothprod763, wboothprod764, wboothprod765, wadd761d, wadd761c );
smul_full_add u501 ( wadd751d, wadd756d, wadd761d, wadd749d, wadd749c );
smul_full_add u502 ( wadd740d, wadd742d, wadd749d, wadd738d, wadd738c );
smul_booth_prod u503 ( x[23], x[24], x[25], y[2], y[3], wboothprod766 );
smul_booth_prod u504 ( x[25], x[26], x[27], y[0], y[1], wboothprod767 );
smul_full_add u505 ( wadd738d, wboothprod766, wboothprod767, wadd736d, wadd736c );
smul_full_add u506 ( wadd684c, wadd732d, wadd736d, wadd730d, wadd730c );
smul_half_add u507 ( wadd682c, wadd730d, wadd728d, wadd728c );
smul_carry_prop u508 ( wadd680d, 1'b0, wcarry769g, wcarry769p );
smul_carry_eval u509 ( wcarry769g, wcarry769p, wcarry721, wcarry768 );
smul_full_add u510 ( wadd680c, wadd728d, wcarry768, wadd726d, wadd726c );
smul_full_add u511 ( wadd740c, wadd742c, wadd749c, wadd779d, wadd779c );
smul_full_add u512 ( wadd734c, wadd738c, wadd779d, wadd777d, wadd777c );
smul_full_add u513 ( wadd732c, wadd736c, wadd777d, wadd775d, wadd775c );
smul_full_add u514 ( wadd744c, wadd751c, wadd756c, wadd785d, wadd785c );
smul_booth_prod u515 ( 1'b0, x[0], x[1], y[27], y[28], wboothprod791 );
smul_booth_prod u516 ( x[1], x[2], x[3], y[25], y[26], wboothprod792 );
smul_booth_prod u517 ( x[3], x[4], x[5], y[23], y[24], wboothprod793 );
smul_full_add u518 ( wboothprod791, wboothprod792, wboothprod793, wadd789d, wadd789c );
smul_booth_prod u519 ( x[5], x[6], x[7], y[21], y[22], wboothprod796 );
smul_booth_prod u520 ( x[7], x[8], x[9], y[19], y[20], wboothprod797 );
smul_booth_prod u521 ( x[9], x[10], x[11], y[17], y[18], wboothprod798 );
smul_full_add u522 ( wboothprod796, wboothprod797, wboothprod798, wadd794d, wadd794c );
smul_full_add u523 ( wadd761c, wadd789d, wadd794d, wadd787d, wadd787c );
smul_booth_prod u524 ( x[11], x[12], x[13], y[15], y[16], wboothprod803 );
smul_booth_prod u525 ( x[13], x[14], x[15], y[13], y[14], wboothprod804 );
smul_booth_prod u526 ( x[15], x[16], x[17], y[11], y[12], wboothprod805 );
smul_full_add u527 ( wboothprod803, wboothprod804, wboothprod805, wadd801d, wadd801c );
smul_booth_prod u528 ( x[17], x[18], x[19], y[9], y[10], wboothprod808 );
smul_booth_prod u529 ( x[19], x[20], x[21], y[7], y[8], wboothprod809 );
smul_booth_prod u530 ( x[21], x[22], x[23], y[5], y[6], wboothprod810 );
smul_full_add u531 ( wboothprod808, wboothprod809, wboothprod810, wadd806d, wadd806c );
smul_booth_prod u532 ( x[23], x[24], x[25], y[3], y[4], wboothprod813 );
smul_booth_prod u533 ( x[25], x[26], x[27], y[1], y[2], wboothprod814 );
smul_booth_prod u534 ( x[27], x[28], x[29], 1'b0, y[0], wboothprod815 );
smul_full_add u535 ( wboothprod813, wboothprod814, wboothprod815, wadd811d, wadd811c );
smul_full_add u536 ( wadd801d, wadd806d, wadd811d, wadd799d, wadd799c );
smul_full_add u537 ( wadd785d, wadd787d, wadd799d, wadd783d, wadd783c );
smul_booth_neg u538 ( x[27], x[28], x[29], wboothneg816 );
smul_half_add u539 ( wadd783d, wboothneg816, wadd781d, wadd781c );
smul_full_add u540 ( wadd730c, wadd775d, wadd781d, wadd773d, wadd773c );
smul_carry_prop u541 ( wadd680c, wadd728d, wcarry822g, wcarry822p );
smul_carry_merge u542 ( wcarry769g, wcarry769p, wcarry822g, wcarry822p, wcarry820g, wcarry820p );
smul_carry_merge u543 ( wcarry722g, wcarry722p, wcarry820g, wcarry820p, wcarry818g, wcarry818p );
smul_carry_eval u544 ( wcarry818g, wcarry818p, wcarry627, wcarry817 );
smul_full_add u545 ( wadd728c, wadd773d, wcarry817, wadd771d, wadd771c );
smul_full_add u546 ( wadd785c, wadd787c, wadd799c, wadd832d, wadd832c );
smul_full_add u547 ( wadd779c, wadd783c, wadd832d, wadd830d, wadd830c );
smul_full_add u548 ( wadd789c, wadd794c, wadd801c, wadd838d, wadd838c );
smul_booth_prod u549 ( 1'b0, x[0], x[1], y[28], y[29], wboothprod844 );
smul_booth_prod u550 ( x[1], x[2], x[3], y[26], y[27], wboothprod845 );
smul_booth_prod u551 ( x[3], x[4], x[5], y[24], y[25], wboothprod846 );
smul_full_add u552 ( wboothprod844, wboothprod845, wboothprod846, wadd842d, wadd842c );
smul_full_add u553 ( wadd806c, wadd811c, wadd842d, wadd840d, wadd840c );
smul_booth_prod u554 ( x[5], x[6], x[7], y[22], y[23], wboothprod851 );
smul_booth_prod u555 ( x[7], x[8], x[9], y[20], y[21], wboothprod852 );
smul_booth_prod u556 ( x[9], x[10], x[11], y[18], y[19], wboothprod853 );
smul_full_add u557 ( wboothprod851, wboothprod852, wboothprod853, wadd849d, wadd849c );
smul_booth_prod u558 ( x[11], x[12], x[13], y[16], y[17], wboothprod856 );
smul_booth_prod u559 ( x[13], x[14], x[15], y[14], y[15], wboothprod857 );
smul_booth_prod u560 ( x[15], x[16], x[17], y[12], y[13], wboothprod858 );
smul_full_add u561 ( wboothprod856, wboothprod857, wboothprod858, wadd854d, wadd854c );
smul_booth_prod u562 ( x[17], x[18], x[19], y[10], y[11], wboothprod861 );
smul_booth_prod u563 ( x[19], x[20], x[21], y[8], y[9], wboothprod862 );
smul_booth_prod u564 ( x[21], x[22], x[23], y[6], y[7], wboothprod863 );
smul_full_add u565 ( wboothprod861, wboothprod862, wboothprod863, wadd859d, wadd859c );
smul_full_add u566 ( wadd849d, wadd854d, wadd859d, wadd847d, wadd847c );
smul_full_add u567 ( wadd838d, wadd840d, wadd847d, wadd836d, wadd836c );
smul_booth_prod u568 ( x[23], x[24], x[25], y[4], y[5], wboothprod866 );
smul_booth_prod u569 ( x[25], x[26], x[27], y[2], y[3], wboothprod867 );
smul_booth_prod u570 ( x[27], x[28], x[29], y[0], y[1], wboothprod868 );
smul_full_add u571 ( wboothprod866, wboothprod867, wboothprod868, wadd864d, wadd864c );
smul_half_add u572 ( wadd836d, wadd864d, wadd834d, wadd834c );
smul_full_add u573 ( wadd777c, wadd830d, wadd834d, wadd828d, wadd828c );
smul_full_add u574 ( wadd775c, wadd781c, wadd828d, wadd826d, wadd826c );
smul_carry_prop u575 ( wadd728c, wadd773d, wcarry870g, wcarry870p );
smul_carry_eval u576 ( wcarry870g, wcarry870p, wcarry817, wcarry869 );
smul_full_add u577 ( wadd773c, wadd826d, wcarry869, wadd824d, wadd824c );
smul_full_add u578 ( wadd838c, wadd840c, wadd847c, wadd880d, wadd880c );
smul_full_add u579 ( wadd832c, wadd836c, wadd880d, wadd878d, wadd878c );
smul_full_add u580 ( wadd830c, wadd834c, wadd878d, wadd876d, wadd876c );
smul_full_add u581 ( wadd842c, wadd849c, wadd854c, wadd886d, wadd886c );
smul_booth_prod u582 ( 1'b0, x[0], x[1], y[29], y[30], wboothprod892 );
smul_booth_prod u583 ( x[1], x[2], x[3], y[27], y[28], wboothprod893 );
smul_booth_prod u584 ( x[3], x[4], x[5], y[25], y[26], wboothprod894 );
smul_full_add u585 ( wboothprod892, wboothprod893, wboothprod894, wadd890d, wadd890c );
smul_full_add u586 ( wadd859c, wadd864c, wadd890d, wadd888d, wadd888c );
smul_booth_prod u587 ( x[5], x[6], x[7], y[23], y[24], wboothprod899 );
smul_booth_prod u588 ( x[7], x[8], x[9], y[21], y[22], wboothprod900 );
smul_booth_prod u589 ( x[9], x[10], x[11], y[19], y[20], wboothprod901 );
smul_full_add u590 ( wboothprod899, wboothprod900, wboothprod901, wadd897d, wadd897c );
smul_booth_prod u591 ( x[11], x[12], x[13], y[17], y[18], wboothprod904 );
smul_booth_prod u592 ( x[13], x[14], x[15], y[15], y[16], wboothprod905 );
smul_booth_prod u593 ( x[15], x[16], x[17], y[13], y[14], wboothprod906 );
smul_full_add u594 ( wboothprod904, wboothprod905, wboothprod906, wadd902d, wadd902c );
smul_booth_prod u595 ( x[17], x[18], x[19], y[11], y[12], wboothprod909 );
smul_booth_prod u596 ( x[19], x[20], x[21], y[9], y[10], wboothprod910 );
smul_booth_prod u597 ( x[21], x[22], x[23], y[7], y[8], wboothprod911 );
smul_full_add u598 ( wboothprod909, wboothprod910, wboothprod911, wadd907d, wadd907c );
smul_full_add u599 ( wadd897d, wadd902d, wadd907d, wadd895d, wadd895c );
smul_full_add u600 ( wadd886d, wadd888d, wadd895d, wadd884d, wadd884c );
smul_booth_prod u601 ( x[23], x[24], x[25], y[5], y[6], wboothprod916 );
smul_booth_prod u602 ( x[25], x[26], x[27], y[3], y[4], wboothprod917 );
smul_booth_prod u603 ( x[27], x[28], x[29], y[1], y[2], wboothprod918 );
smul_full_add u604 ( wboothprod916, wboothprod917, wboothprod918, wadd914d, wadd914c );
smul_booth_prod u605 ( x[29], x[30], x[31], 1'b0, y[0], wboothprod919 );
smul_booth_neg u606 ( x[29], x[30], x[31], wboothneg920 );
smul_full_add u607 ( wadd914d, wboothprod919, wboothneg920, wadd912d, wadd912c );
smul_half_add u608 ( wadd884d, wadd912d, wadd882d, wadd882c );
smul_full_add u609 ( wadd828c, wadd876d, wadd882d, wadd874d, wadd874c );
smul_carry_prop u610 ( wadd773c, wadd826d, wcarry924g, wcarry924p );
smul_carry_merge u611 ( wcarry870g, wcarry870p, wcarry924g, wcarry924p, wcarry922g, wcarry922p );
smul_carry_eval u612 ( wcarry922g, wcarry922p, wcarry817, wcarry921 );
smul_full_add u613 ( wadd826c, wadd874d, wcarry921, wadd872d, wadd872c );
smul_full_add u614 ( wadd886c, wadd888c, wadd895c, wadd934d, wadd934c );
smul_full_add u615 ( wadd880c, wadd884c, wadd934d, wadd932d, wadd932c );
smul_full_add u616 ( wadd890c, wadd897c, wadd902c, wadd940d, wadd940c );
smul_booth_prod u617 ( 1'b0, x[0], x[1], y[30], y[31], wboothprod946 );
smul_booth_prod u618 ( x[1], x[2], x[3], y[28], y[29], wboothprod947 );
smul_booth_prod u619 ( x[3], x[4], x[5], y[26], y[27], wboothprod948 );
smul_full_add u620 ( wboothprod946, wboothprod947, wboothprod948, wadd944d, wadd944c );
smul_full_add u621 ( wadd907c, wadd914c, wadd944d, wadd942d, wadd942c );
smul_full_add u622 ( wadd912c, wadd940d, wadd942d, wadd938d, wadd938c );
smul_booth_prod u623 ( x[5], x[6], x[7], y[24], y[25], wboothprod955 );
smul_booth_prod u624 ( x[7], x[8], x[9], y[22], y[23], wboothprod956 );
smul_booth_prod u625 ( x[9], x[10], x[11], y[20], y[21], wboothprod957 );
smul_full_add u626 ( wboothprod955, wboothprod956, wboothprod957, wadd953d, wadd953c );
smul_booth_prod u627 ( x[11], x[12], x[13], y[18], y[19], wboothprod960 );
smul_booth_prod u628 ( x[13], x[14], x[15], y[16], y[17], wboothprod961 );
smul_booth_prod u629 ( x[15], x[16], x[17], y[14], y[15], wboothprod962 );
smul_full_add u630 ( wboothprod960, wboothprod961, wboothprod962, wadd958d, wadd958c );
smul_booth_prod u631 ( x[17], x[18], x[19], y[12], y[13], wboothprod965 );
smul_booth_prod u632 ( x[19], x[20], x[21], y[10], y[11], wboothprod966 );
smul_booth_prod u633 ( x[21], x[22], x[23], y[8], y[9], wboothprod967 );
smul_full_add u634 ( wboothprod965, wboothprod966, wboothprod967, wadd963d, wadd963c );
smul_full_add u635 ( wadd953d, wadd958d, wadd963d, wadd951d, wadd951c );
smul_booth_prod u636 ( x[23], x[24], x[25], y[6], y[7], wboothprod970 );
smul_booth_prod u637 ( x[25], x[26], x[27], y[4], y[5], wboothprod971 );
smul_booth_prod u638 ( x[27], x[28], x[29], y[2], y[3], wboothprod972 );
smul_full_add u639 ( wboothprod970, wboothprod971, wboothprod972, wadd968d, wadd968c );
smul_booth_prod u640 ( x[29], x[30], x[31], y[0], y[1], wboothprod973 );
smul_full_add u641 ( wadd951d, wadd968d, wboothprod973, wadd949d, wadd949c );
smul_half_add u642 ( wadd938d, wadd949d, wadd936d, wadd936c );
smul_full_add u643 ( wadd878c, wadd932d, wadd936d, wadd930d, wadd930c );
smul_full_add u644 ( wadd876c, wadd882c, wadd930d, wadd928d, wadd928c );
smul_carry_prop u645 ( wadd826c, wadd874d, wcarry975g, wcarry975p );
smul_carry_eval u646 ( wcarry975g, wcarry975p, wcarry921, wcarry974 );
smul_full_add u647 ( wadd874c, wadd928d, wcarry974, wadd926d, wadd926c );
smul_full_add u648 ( wadd934c, wadd938c, wadd949c, wadd983d, wadd983c );
smul_full_add u649 ( wadd932c, wadd936c, wadd983d, wadd981d, wadd981c );
smul_full_add u650 ( wadd940c, wadd942c, wadd951c, wadd987d, wadd987c );
smul_full_add u651 ( wadd944c, wadd953c, wadd958c, wadd991d, wadd991c );
smul_booth_prod u652 ( 1'b0, x[0], x[1], y[31], y[31], wboothprod997 );
smul_booth_prod u653 ( x[1], x[2], x[3], y[29], y[30], wboothprod998 );
smul_booth_prod u654 ( x[3], x[4], x[5], y[27], y[28], wboothprod999 );
smul_full_add u655 ( wboothprod997, wboothprod998, wboothprod999, wadd995d, wadd995c );
smul_full_add u656 ( wadd963c, wadd968c, wadd995d, wadd993d, wadd993c );
smul_booth_prod u657 ( x[5], x[6], x[7], y[25], y[26], wboothprod1004 );
smul_booth_prod u658 ( x[7], x[8], x[9], y[23], y[24], wboothprod1005 );
smul_booth_prod u659 ( x[9], x[10], x[11], y[21], y[22], wboothprod1006 );
smul_full_add u660 ( wboothprod1004, wboothprod1005, wboothprod1006, wadd1002d, wadd1002c );
smul_booth_prod u661 ( x[11], x[12], x[13], y[19], y[20], wboothprod1009 );
smul_booth_prod u662 ( x[13], x[14], x[15], y[17], y[18], wboothprod1010 );
smul_booth_prod u663 ( x[15], x[16], x[17], y[15], y[16], wboothprod1011 );
smul_full_add u664 ( wboothprod1009, wboothprod1010, wboothprod1011, wadd1007d, wadd1007c );
smul_booth_prod u665 ( x[17], x[18], x[19], y[13], y[14], wboothprod1014 );
smul_booth_prod u666 ( x[19], x[20], x[21], y[11], y[12], wboothprod1015 );
smul_booth_prod u667 ( x[21], x[22], x[23], y[9], y[10], wboothprod1016 );
smul_full_add u668 ( wboothprod1014, wboothprod1015, wboothprod1016, wadd1012d, wadd1012c );
smul_full_add u669 ( wadd1002d, wadd1007d, wadd1012d, wadd1000d, wadd1000c );
smul_full_add u670 ( wadd991d, wadd993d, wadd1000d, wadd989d, wadd989c );
smul_booth_prod u671 ( x[23], x[24], x[25], y[7], y[8], wboothprod1021 );
smul_booth_prod u672 ( x[25], x[26], x[27], y[5], y[6], wboothprod1022 );
smul_booth_prod u673 ( x[27], x[28], x[29], y[3], y[4], wboothprod1023 );
smul_full_add u674 ( wboothprod1021, wboothprod1022, wboothprod1023, wadd1019d, wadd1019c );
smul_booth_prod u675 ( x[29], x[30], x[31], y[1], y[2], wboothprod1024 );
smul_half_add u676 ( wadd1019d, wboothprod1024, wadd1017d, wadd1017c );
smul_full_add u677 ( wadd987d, wadd989d, wadd1017d, wadd985d, wadd985c );
smul_full_add u678 ( wadd930c, wadd981d, wadd985d, wadd979d, wadd979c );
smul_carry_prop u679 ( wadd874c, wadd928d, wcarry1036g, wcarry1036p );
smul_carry_merge u680 ( wcarry975g, wcarry975p, wcarry1036g, wcarry1036p, wcarry1034g, wcarry1034p );
smul_carry_merge u681 ( wcarry922g, wcarry922p, wcarry1034g, wcarry1034p, wcarry1032g, wcarry1032p );
smul_carry_merge u682 ( wcarry818g, wcarry818p, wcarry1032g, wcarry1032p, wcarry1030g, wcarry1030p );
smul_carry_merge u683 ( wcarry628g, wcarry628p, wcarry1030g, wcarry1030p, wcarry1028g, wcarry1028p );
smul_carry_merge u684 ( wcarry320g, wcarry320p, wcarry1028g, wcarry1028p, wcarry1026g, wcarry1026p );
smul_carry_eval u685 ( wcarry1026g, wcarry1026p, 1'b0, wcarry1025 );
smul_full_add u686 ( wadd928c, wadd979d, wcarry1025, wadd977d, wadd977c );
smul_full_add u687 ( wadd987c, wadd989c, wadd1017c, wadd1044d, wadd1044c );
smul_full_add u688 ( wadd983c, wadd985c, wadd1044d, wadd1042d, wadd1042c );
smul_full_add u689 ( wadd991c, wadd993c, wadd1000c, wadd1048d, wadd1048c );
smul_full_add u690 ( wadd995c, wadd1002c, wadd1007c, wadd1052d, wadd1052c );
smul_booth_prod u691 ( x[1], x[2], x[3], y[30], y[31], wboothprod1058 );
smul_booth_prod u692 ( x[3], x[4], x[5], y[28], y[29], wboothprod1059 );
smul_full_add u693 ( wboothprod997, wboothprod1058, wboothprod1059, wadd1056d, wadd1056c );
smul_full_add u694 ( wadd1012c, wadd1019c, wadd1056d, wadd1054d, wadd1054c );
smul_booth_prod u695 ( x[5], x[6], x[7], y[26], y[27], wboothprod1064 );
smul_booth_prod u696 ( x[7], x[8], x[9], y[24], y[25], wboothprod1065 );
smul_booth_prod u697 ( x[9], x[10], x[11], y[22], y[23], wboothprod1066 );
smul_full_add u698 ( wboothprod1064, wboothprod1065, wboothprod1066, wadd1062d, wadd1062c );
smul_booth_prod u699 ( x[11], x[12], x[13], y[20], y[21], wboothprod1069 );
smul_booth_prod u700 ( x[13], x[14], x[15], y[18], y[19], wboothprod1070 );
smul_booth_prod u701 ( x[15], x[16], x[17], y[16], y[17], wboothprod1071 );
smul_full_add u702 ( wboothprod1069, wboothprod1070, wboothprod1071, wadd1067d, wadd1067c );
smul_booth_prod u703 ( x[17], x[18], x[19], y[14], y[15], wboothprod1074 );
smul_booth_prod u704 ( x[19], x[20], x[21], y[12], y[13], wboothprod1075 );
smul_booth_prod u705 ( x[21], x[22], x[23], y[10], y[11], wboothprod1076 );
smul_full_add u706 ( wboothprod1074, wboothprod1075, wboothprod1076, wadd1072d, wadd1072c );
smul_full_add u707 ( wadd1062d, wadd1067d, wadd1072d, wadd1060d, wadd1060c );
smul_full_add u708 ( wadd1052d, wadd1054d, wadd1060d, wadd1050d, wadd1050c );
smul_booth_prod u709 ( x[23], x[24], x[25], y[8], y[9], wboothprod1081 );
smul_booth_prod u710 ( x[25], x[26], x[27], y[6], y[7], wboothprod1082 );
smul_booth_prod u711 ( x[27], x[28], x[29], y[4], y[5], wboothprod1083 );
smul_full_add u712 ( wboothprod1081, wboothprod1082, wboothprod1083, wadd1079d, wadd1079c );
smul_booth_prod u713 ( x[29], x[30], x[31], y[2], y[3], wboothprod1084 );
smul_half_add u714 ( wadd1079d, wboothprod1084, wadd1077d, wadd1077c );
smul_full_add u715 ( wadd1048d, wadd1050d, wadd1077d, wadd1046d, wadd1046c );
smul_full_add u716 ( wadd981c, wadd1042d, wadd1046d, wadd1040d, wadd1040c );
smul_carry_prop u717 ( wadd928c, wadd979d, wcarry1086g, wcarry1086p );
smul_carry_eval u718 ( wcarry1086g, wcarry1086p, wcarry1025, wcarry1085 );
smul_full_add u719 ( wadd979c, wadd1040d, wcarry1085, wadd1038d, wadd1038c );
smul_full_add u720 ( wadd1048c, wadd1050c, wadd1077c, wadd1094d, wadd1094c );
smul_full_add u721 ( wadd1044c, wadd1046c, wadd1094d, wadd1092d, wadd1092c );
smul_full_add u722 ( wadd1052c, wadd1054c, wadd1060c, wadd1098d, wadd1098c );
smul_full_add u723 ( wadd1056c, wadd1062c, wadd1067c, wadd1102d, wadd1102c );
smul_inverter u724 ( wboothprod997, winv1108 );
smul_booth_prod u725 ( x[1], x[2], x[3], y[31], y[31], wboothprod1110 );
smul_inverter u726 ( wboothprod1110, winv1109 );
smul_booth_prod u727 ( x[3], x[4], x[5], y[29], y[30], wboothprod1111 );
smul_full_add u728 ( winv1108, winv1109, wboothprod1111, wadd1106d, wadd1106c );
smul_full_add u729 ( wadd1072c, wadd1079c, wadd1106d, wadd1104d, wadd1104c );
smul_booth_prod u730 ( x[5], x[6], x[7], y[27], y[28], wboothprod1116 );
smul_booth_prod u731 ( x[7], x[8], x[9], y[25], y[26], wboothprod1117 );
smul_booth_prod u732 ( x[9], x[10], x[11], y[23], y[24], wboothprod1118 );
smul_full_add u733 ( wboothprod1116, wboothprod1117, wboothprod1118, wadd1114d, wadd1114c );
smul_booth_prod u734 ( x[11], x[12], x[13], y[21], y[22], wboothprod1121 );
smul_booth_prod u735 ( x[13], x[14], x[15], y[19], y[20], wboothprod1122 );
smul_booth_prod u736 ( x[15], x[16], x[17], y[17], y[18], wboothprod1123 );
smul_full_add u737 ( wboothprod1121, wboothprod1122, wboothprod1123, wadd1119d, wadd1119c );
smul_booth_prod u738 ( x[17], x[18], x[19], y[15], y[16], wboothprod1126 );
smul_booth_prod u739 ( x[19], x[20], x[21], y[13], y[14], wboothprod1127 );
smul_booth_prod u740 ( x[21], x[22], x[23], y[11], y[12], wboothprod1128 );
smul_full_add u741 ( wboothprod1126, wboothprod1127, wboothprod1128, wadd1124d, wadd1124c );
smul_full_add u742 ( wadd1114d, wadd1119d, wadd1124d, wadd1112d, wadd1112c );
smul_full_add u743 ( wadd1102d, wadd1104d, wadd1112d, wadd1100d, wadd1100c );
smul_booth_prod u744 ( x[23], x[24], x[25], y[9], y[10], wboothprod1133 );
smul_booth_prod u745 ( x[25], x[26], x[27], y[7], y[8], wboothprod1134 );
smul_booth_prod u746 ( x[27], x[28], x[29], y[5], y[6], wboothprod1135 );
smul_full_add u747 ( wboothprod1133, wboothprod1134, wboothprod1135, wadd1131d, wadd1131c );
smul_booth_prod u748 ( x[29], x[30], x[31], y[3], y[4], wboothprod1136 );
smul_half_add u749 ( wadd1131d, wboothprod1136, wadd1129d, wadd1129c );
smul_full_add u750 ( wadd1098d, wadd1100d, wadd1129d, wadd1096d, wadd1096c );
smul_full_add u751 ( wadd1042c, wadd1092d, wadd1096d, wadd1090d, wadd1090c );
smul_carry_prop u752 ( wadd979c, wadd1040d, wcarry1140g, wcarry1140p );
smul_carry_merge u753 ( wcarry1086g, wcarry1086p, wcarry1140g, wcarry1140p, wcarry1138g, wcarry1138p );
smul_carry_eval u754 ( wcarry1138g, wcarry1138p, wcarry1025, wcarry1137 );
smul_full_add u755 ( wadd1040c, wadd1090d, wcarry1137, wadd1088d, wadd1088c );
smul_full_add u756 ( wadd1098c, wadd1100c, wadd1129c, wadd1148d, wadd1148c );
smul_full_add u757 ( wadd1094c, wadd1096c, wadd1148d, wadd1146d, wadd1146c );
smul_full_add u758 ( wadd1102c, wadd1104c, wadd1112c, wadd1152d, wadd1152c );
smul_full_add u759 ( wadd1106c, wadd1114c, wadd1119c, wadd1156d, wadd1156c );
smul_booth_prod u760 ( x[3], x[4], x[5], y[30], y[31], wboothprod1162 );
smul_booth_prod u761 ( x[5], x[6], x[7], y[28], y[29], wboothprod1163 );
smul_full_add u762 ( 1'b1, wboothprod1162, wboothprod1163, wadd1160d, wadd1160c );
smul_full_add u763 ( wadd1124c, wadd1131c, wadd1160d, wadd1158d, wadd1158c );
smul_booth_prod u764 ( x[7], x[8], x[9], y[26], y[27], wboothprod1168 );
smul_booth_prod u765 ( x[9], x[10], x[11], y[24], y[25], wboothprod1169 );
smul_booth_prod u766 ( x[11], x[12], x[13], y[22], y[23], wboothprod1170 );
smul_full_add u767 ( wboothprod1168, wboothprod1169, wboothprod1170, wadd1166d, wadd1166c );
smul_booth_prod u768 ( x[13], x[14], x[15], y[20], y[21], wboothprod1173 );
smul_booth_prod u769 ( x[15], x[16], x[17], y[18], y[19], wboothprod1174 );
smul_booth_prod u770 ( x[17], x[18], x[19], y[16], y[17], wboothprod1175 );
smul_full_add u771 ( wboothprod1173, wboothprod1174, wboothprod1175, wadd1171d, wadd1171c );
smul_booth_prod u772 ( x[19], x[20], x[21], y[14], y[15], wboothprod1178 );
smul_booth_prod u773 ( x[21], x[22], x[23], y[12], y[13], wboothprod1179 );
smul_booth_prod u774 ( x[23], x[24], x[25], y[10], y[11], wboothprod1180 );
smul_full_add u775 ( wboothprod1178, wboothprod1179, wboothprod1180, wadd1176d, wadd1176c );
smul_full_add u776 ( wadd1166d, wadd1171d, wadd1176d, wadd1164d, wadd1164c );
smul_full_add u777 ( wadd1156d, wadd1158d, wadd1164d, wadd1154d, wadd1154c );
smul_booth_prod u778 ( x[25], x[26], x[27], y[8], y[9], wboothprod1183 );
smul_booth_prod u779 ( x[27], x[28], x[29], y[6], y[7], wboothprod1184 );
smul_booth_prod u780 ( x[29], x[30], x[31], y[4], y[5], wboothprod1185 );
smul_full_add u781 ( wboothprod1183, wboothprod1184, wboothprod1185, wadd1181d, wadd1181c );
smul_full_add u782 ( wadd1152d, wadd1154d, wadd1181d, wadd1150d, wadd1150c );
smul_full_add u783 ( wadd1092c, wadd1146d, wadd1150d, wadd1144d, wadd1144c );
smul_carry_prop u784 ( wadd1040c, wadd1090d, wcarry1187g, wcarry1187p );
smul_carry_eval u785 ( wcarry1187g, wcarry1187p, wcarry1137, wcarry1186 );
smul_full_add u786 ( wadd1090c, wadd1144d, wcarry1186, wadd1142d, wadd1142c );
smul_full_add u787 ( wadd1156c, wadd1158c, wadd1164c, wadd1197d, wadd1197c );
smul_full_add u788 ( wadd1152c, wadd1154c, wadd1197d, wadd1195d, wadd1195c );
smul_full_add u789 ( wadd1148c, wadd1150c, wadd1195d, wadd1193d, wadd1193c );
smul_full_add u790 ( wadd1160c, wadd1166c, wadd1171c, wadd1203d, wadd1203c );
smul_booth_prod u791 ( x[3], x[4], x[5], y[31], y[31], wboothprod1210 );
smul_inverter u792 ( wboothprod1210, winv1209 );
smul_booth_prod u793 ( x[5], x[6], x[7], y[29], y[30], wboothprod1211 );
smul_booth_prod u794 ( x[7], x[8], x[9], y[27], y[28], wboothprod1212 );
smul_full_add u795 ( winv1209, wboothprod1211, wboothprod1212, wadd1207d, wadd1207c );
smul_full_add u796 ( wadd1176c, wadd1181c, wadd1207d, wadd1205d, wadd1205c );
smul_booth_prod u797 ( x[9], x[10], x[11], y[25], y[26], wboothprod1217 );
smul_booth_prod u798 ( x[11], x[12], x[13], y[23], y[24], wboothprod1218 );
smul_booth_prod u799 ( x[13], x[14], x[15], y[21], y[22], wboothprod1219 );
smul_full_add u800 ( wboothprod1217, wboothprod1218, wboothprod1219, wadd1215d, wadd1215c );
smul_booth_prod u801 ( x[15], x[16], x[17], y[19], y[20], wboothprod1222 );
smul_booth_prod u802 ( x[17], x[18], x[19], y[17], y[18], wboothprod1223 );
smul_booth_prod u803 ( x[19], x[20], x[21], y[15], y[16], wboothprod1224 );
smul_full_add u804 ( wboothprod1222, wboothprod1223, wboothprod1224, wadd1220d, wadd1220c );
smul_booth_prod u805 ( x[21], x[22], x[23], y[13], y[14], wboothprod1227 );
smul_booth_prod u806 ( x[23], x[24], x[25], y[11], y[12], wboothprod1228 );
smul_booth_prod u807 ( x[25], x[26], x[27], y[9], y[10], wboothprod1229 );
smul_full_add u808 ( wboothprod1227, wboothprod1228, wboothprod1229, wadd1225d, wadd1225c );
smul_full_add u809 ( wadd1215d, wadd1220d, wadd1225d, wadd1213d, wadd1213c );
smul_full_add u810 ( wadd1203d, wadd1205d, wadd1213d, wadd1201d, wadd1201c );
smul_booth_prod u811 ( x[27], x[28], x[29], y[7], y[8], wboothprod1230 );
smul_booth_prod u812 ( x[29], x[30], x[31], y[5], y[6], wboothprod1231 );
smul_full_add u813 ( wadd1201d, wboothprod1230, wboothprod1231, wadd1199d, wadd1199c );
smul_full_add u814 ( wadd1146c, wadd1193d, wadd1199d, wadd1191d, wadd1191c );
smul_carry_prop u815 ( wadd1090c, wadd1144d, wcarry1237g, wcarry1237p );
smul_carry_merge u816 ( wcarry1187g, wcarry1187p, wcarry1237g, wcarry1237p, wcarry1235g, wcarry1235p );
smul_carry_merge u817 ( wcarry1138g, wcarry1138p, wcarry1235g, wcarry1235p, wcarry1233g, wcarry1233p );
smul_carry_eval u818 ( wcarry1233g, wcarry1233p, wcarry1025, wcarry1232 );
smul_full_add u819 ( wadd1144c, wadd1191d, wcarry1232, wadd1189d, wadd1189c );
smul_full_add u820 ( wadd1203c, wadd1205c, wadd1213c, wadd1247d, wadd1247c );
smul_full_add u821 ( wadd1197c, wadd1201c, wadd1247d, wadd1245d, wadd1245c );
smul_full_add u822 ( wadd1195c, wadd1199c, wadd1245d, wadd1243d, wadd1243c );
smul_full_add u823 ( wadd1207c, wadd1215c, wadd1220c, wadd1251d, wadd1251c );
smul_booth_prod u824 ( x[5], x[6], x[7], y[30], y[31], wboothprod1257 );
smul_booth_prod u825 ( x[7], x[8], x[9], y[28], y[29], wboothprod1258 );
smul_full_add u826 ( 1'b1, wboothprod1257, wboothprod1258, wadd1255d, wadd1255c );
smul_booth_prod u827 ( x[9], x[10], x[11], y[26], y[27], wboothprod1261 );
smul_booth_prod u828 ( x[11], x[12], x[13], y[24], y[25], wboothprod1262 );
smul_booth_prod u829 ( x[13], x[14], x[15], y[22], y[23], wboothprod1263 );
smul_full_add u830 ( wboothprod1261, wboothprod1262, wboothprod1263, wadd1259d, wadd1259c );
smul_full_add u831 ( wadd1225c, wadd1255d, wadd1259d, wadd1253d, wadd1253c );
smul_booth_prod u832 ( x[15], x[16], x[17], y[20], y[21], wboothprod1268 );
smul_booth_prod u833 ( x[17], x[18], x[19], y[18], y[19], wboothprod1269 );
smul_booth_prod u834 ( x[19], x[20], x[21], y[16], y[17], wboothprod1270 );
smul_full_add u835 ( wboothprod1268, wboothprod1269, wboothprod1270, wadd1266d, wadd1266c );
smul_booth_prod u836 ( x[21], x[22], x[23], y[14], y[15], wboothprod1273 );
smul_booth_prod u837 ( x[23], x[24], x[25], y[12], y[13], wboothprod1274 );
smul_booth_prod u838 ( x[25], x[26], x[27], y[10], y[11], wboothprod1275 );
smul_full_add u839 ( wboothprod1273, wboothprod1274, wboothprod1275, wadd1271d, wadd1271c );
smul_booth_prod u840 ( x[27], x[28], x[29], y[8], y[9], wboothprod1278 );
smul_booth_prod u841 ( x[29], x[30], x[31], y[6], y[7], wboothprod1279 );
smul_half_add u842 ( wboothprod1278, wboothprod1279, wadd1276d, wadd1276c );
smul_full_add u843 ( wadd1266d, wadd1271d, wadd1276d, wadd1264d, wadd1264c );
smul_full_add u844 ( wadd1251d, wadd1253d, wadd1264d, wadd1249d, wadd1249c );
smul_full_add u845 ( wadd1193c, wadd1243d, wadd1249d, wadd1241d, wadd1241c );
smul_carry_prop u846 ( wadd1144c, wadd1191d, wcarry1281g, wcarry1281p );
smul_carry_eval u847 ( wcarry1281g, wcarry1281p, wcarry1232, wcarry1280 );
smul_full_add u848 ( wadd1191c, wadd1241d, wcarry1280, wadd1239d, wadd1239c );
smul_full_add u849 ( wadd1251c, wadd1253c, wadd1264c, wadd1291d, wadd1291c );
smul_full_add u850 ( wadd1247c, wadd1249c, wadd1291d, wadd1289d, wadd1289c );
smul_full_add u851 ( wadd1255c, wadd1259c, wadd1266c, wadd1297d, wadd1297c );
smul_booth_prod u852 ( x[5], x[6], x[7], y[31], y[31], wboothprod1304 );
smul_inverter u853 ( wboothprod1304, winv1303 );
smul_booth_prod u854 ( x[7], x[8], x[9], y[29], y[30], wboothprod1305 );
smul_booth_prod u855 ( x[9], x[10], x[11], y[27], y[28], wboothprod1306 );
smul_full_add u856 ( winv1303, wboothprod1305, wboothprod1306, wadd1301d, wadd1301c );
smul_full_add u857 ( wadd1271c, wadd1276c, wadd1301d, wadd1299d, wadd1299c );
smul_booth_prod u858 ( x[11], x[12], x[13], y[25], y[26], wboothprod1311 );
smul_booth_prod u859 ( x[13], x[14], x[15], y[23], y[24], wboothprod1312 );
smul_booth_prod u860 ( x[15], x[16], x[17], y[21], y[22], wboothprod1313 );
smul_full_add u861 ( wboothprod1311, wboothprod1312, wboothprod1313, wadd1309d, wadd1309c );
smul_booth_prod u862 ( x[17], x[18], x[19], y[19], y[20], wboothprod1316 );
smul_booth_prod u863 ( x[19], x[20], x[21], y[17], y[18], wboothprod1317 );
smul_booth_prod u864 ( x[21], x[22], x[23], y[15], y[16], wboothprod1318 );
smul_full_add u865 ( wboothprod1316, wboothprod1317, wboothprod1318, wadd1314d, wadd1314c );
smul_booth_prod u866 ( x[23], x[24], x[25], y[13], y[14], wboothprod1321 );
smul_booth_prod u867 ( x[25], x[26], x[27], y[11], y[12], wboothprod1322 );
smul_booth_prod u868 ( x[27], x[28], x[29], y[9], y[10], wboothprod1323 );
smul_full_add u869 ( wboothprod1321, wboothprod1322, wboothprod1323, wadd1319d, wadd1319c );
smul_full_add u870 ( wadd1309d, wadd1314d, wadd1319d, wadd1307d, wadd1307c );
smul_full_add u871 ( wadd1297d, wadd1299d, wadd1307d, wadd1295d, wadd1295c );
smul_booth_prod u872 ( x[29], x[30], x[31], y[7], y[8], wboothprod1324 );
smul_half_add u873 ( wadd1295d, wboothprod1324, wadd1293d, wadd1293c );
smul_full_add u874 ( wadd1245c, wadd1289d, wadd1293d, wadd1287d, wadd1287c );
smul_half_add u875 ( wadd1243c, wadd1287d, wadd1285d, wadd1285c );
smul_carry_prop u876 ( wadd1191c, wadd1241d, wcarry1328g, wcarry1328p );
smul_carry_merge u877 ( wcarry1281g, wcarry1281p, wcarry1328g, wcarry1328p, wcarry1326g, wcarry1326p );
smul_carry_eval u878 ( wcarry1326g, wcarry1326p, wcarry1232, wcarry1325 );
smul_full_add u879 ( wadd1241c, wadd1285d, wcarry1325, wadd1283d, wadd1283c );
smul_full_add u880 ( wadd1297c, wadd1299c, wadd1307c, wadd1338d, wadd1338c );
smul_full_add u881 ( wadd1291c, wadd1295c, wadd1338d, wadd1336d, wadd1336c );
smul_full_add u882 ( wadd1289c, wadd1293c, wadd1336d, wadd1334d, wadd1334c );
smul_full_add u883 ( wadd1301c, wadd1309c, wadd1314c, wadd1342d, wadd1342c );
smul_booth_prod u884 ( x[7], x[8], x[9], y[30], y[31], wboothprod1348 );
smul_booth_prod u885 ( x[9], x[10], x[11], y[28], y[29], wboothprod1349 );
smul_full_add u886 ( 1'b1, wboothprod1348, wboothprod1349, wadd1346d, wadd1346c );
smul_booth_prod u887 ( x[11], x[12], x[13], y[26], y[27], wboothprod1352 );
smul_booth_prod u888 ( x[13], x[14], x[15], y[24], y[25], wboothprod1353 );
smul_booth_prod u889 ( x[15], x[16], x[17], y[22], y[23], wboothprod1354 );
smul_full_add u890 ( wboothprod1352, wboothprod1353, wboothprod1354, wadd1350d, wadd1350c );
smul_full_add u891 ( wadd1319c, wadd1346d, wadd1350d, wadd1344d, wadd1344c );
smul_booth_prod u892 ( x[17], x[18], x[19], y[20], y[21], wboothprod1359 );
smul_booth_prod u893 ( x[19], x[20], x[21], y[18], y[19], wboothprod1360 );
smul_booth_prod u894 ( x[21], x[22], x[23], y[16], y[17], wboothprod1361 );
smul_full_add u895 ( wboothprod1359, wboothprod1360, wboothprod1361, wadd1357d, wadd1357c );
smul_booth_prod u896 ( x[23], x[24], x[25], y[14], y[15], wboothprod1364 );
smul_booth_prod u897 ( x[25], x[26], x[27], y[12], y[13], wboothprod1365 );
smul_booth_prod u898 ( x[27], x[28], x[29], y[10], y[11], wboothprod1366 );
smul_full_add u899 ( wboothprod1364, wboothprod1365, wboothprod1366, wadd1362d, wadd1362c );
smul_booth_prod u900 ( x[29], x[30], x[31], y[8], y[9], wboothprod1367 );
smul_full_add u901 ( wadd1357d, wadd1362d, wboothprod1367, wadd1355d, wadd1355c );
smul_full_add u902 ( wadd1342d, wadd1344d, wadd1355d, wadd1340d, wadd1340c );
smul_full_add u903 ( wadd1287c, wadd1334d, wadd1340d, wadd1332d, wadd1332c );
smul_carry_prop u904 ( wadd1241c, wadd1285d, wcarry1369g, wcarry1369p );
smul_carry_eval u905 ( wcarry1369g, wcarry1369p, wcarry1325, wcarry1368 );
smul_full_add u906 ( wadd1285c, wadd1332d, wcarry1368, wadd1330d, wadd1330c );
smul_full_add u907 ( wadd1342c, wadd1344c, wadd1355c, wadd1379d, wadd1379c );
smul_full_add u908 ( wadd1338c, wadd1340c, wadd1379d, wadd1377d, wadd1377c );
smul_full_add u909 ( wadd1346c, wadd1350c, wadd1357c, wadd1383d, wadd1383c );
smul_booth_prod u910 ( x[7], x[8], x[9], y[31], y[31], wboothprod1390 );
smul_inverter u911 ( wboothprod1390, winv1389 );
smul_booth_prod u912 ( x[9], x[10], x[11], y[29], y[30], wboothprod1391 );
smul_booth_prod u913 ( x[11], x[12], x[13], y[27], y[28], wboothprod1392 );
smul_full_add u914 ( winv1389, wboothprod1391, wboothprod1392, wadd1387d, wadd1387c );
smul_booth_prod u915 ( x[13], x[14], x[15], y[25], y[26], wboothprod1395 );
smul_booth_prod u916 ( x[15], x[16], x[17], y[23], y[24], wboothprod1396 );
smul_booth_prod u917 ( x[17], x[18], x[19], y[21], y[22], wboothprod1397 );
smul_full_add u918 ( wboothprod1395, wboothprod1396, wboothprod1397, wadd1393d, wadd1393c );
smul_full_add u919 ( wadd1362c, wadd1387d, wadd1393d, wadd1385d, wadd1385c );
smul_booth_prod u920 ( x[19], x[20], x[21], y[19], y[20], wboothprod1402 );
smul_booth_prod u921 ( x[21], x[22], x[23], y[17], y[18], wboothprod1403 );
smul_booth_prod u922 ( x[23], x[24], x[25], y[15], y[16], wboothprod1404 );
smul_full_add u923 ( wboothprod1402, wboothprod1403, wboothprod1404, wadd1400d, wadd1400c );
smul_booth_prod u924 ( x[25], x[26], x[27], y[13], y[14], wboothprod1407 );
smul_booth_prod u925 ( x[27], x[28], x[29], y[11], y[12], wboothprod1408 );
smul_booth_prod u926 ( x[29], x[30], x[31], y[9], y[10], wboothprod1409 );
smul_full_add u927 ( wboothprod1407, wboothprod1408, wboothprod1409, wadd1405d, wadd1405c );
smul_half_add u928 ( wadd1400d, wadd1405d, wadd1398d, wadd1398c );
smul_full_add u929 ( wadd1383d, wadd1385d, wadd1398d, wadd1381d, wadd1381c );
smul_full_add u930 ( wadd1336c, wadd1377d, wadd1381d, wadd1375d, wadd1375c );
smul_half_add u931 ( wadd1334c, wadd1375d, wadd1373d, wadd1373c );
smul_carry_prop u932 ( wadd1285c, wadd1332d, wcarry1417g, wcarry1417p );
smul_carry_merge u933 ( wcarry1369g, wcarry1369p, wcarry1417g, wcarry1417p, wcarry1415g, wcarry1415p );
smul_carry_merge u934 ( wcarry1326g, wcarry1326p, wcarry1415g, wcarry1415p, wcarry1413g, wcarry1413p );
smul_carry_merge u935 ( wcarry1233g, wcarry1233p, wcarry1413g, wcarry1413p, wcarry1411g, wcarry1411p );
smul_carry_eval u936 ( wcarry1411g, wcarry1411p, wcarry1025, wcarry1410 );
smul_full_add u937 ( wadd1332c, wadd1373d, wcarry1410, wadd1371d, wadd1371c );
smul_full_add u938 ( wadd1383c, wadd1385c, wadd1398c, wadd1427d, wadd1427c );
smul_full_add u939 ( wadd1379c, wadd1381c, wadd1427d, wadd1425d, wadd1425c );
smul_full_add u940 ( wadd1387c, wadd1393c, wadd1400c, wadd1431d, wadd1431c );
smul_booth_prod u941 ( x[9], x[10], x[11], y[30], y[31], wboothprod1437 );
smul_booth_prod u942 ( x[11], x[12], x[13], y[28], y[29], wboothprod1438 );
smul_full_add u943 ( 1'b1, wboothprod1437, wboothprod1438, wadd1435d, wadd1435c );
smul_booth_prod u944 ( x[13], x[14], x[15], y[26], y[27], wboothprod1441 );
smul_booth_prod u945 ( x[15], x[16], x[17], y[24], y[25], wboothprod1442 );
smul_booth_prod u946 ( x[17], x[18], x[19], y[22], y[23], wboothprod1443 );
smul_full_add u947 ( wboothprod1441, wboothprod1442, wboothprod1443, wadd1439d, wadd1439c );
smul_full_add u948 ( wadd1405c, wadd1435d, wadd1439d, wadd1433d, wadd1433c );
smul_booth_prod u949 ( x[19], x[20], x[21], y[20], y[21], wboothprod1448 );
smul_booth_prod u950 ( x[21], x[22], x[23], y[18], y[19], wboothprod1449 );
smul_booth_prod u951 ( x[23], x[24], x[25], y[16], y[17], wboothprod1450 );
smul_full_add u952 ( wboothprod1448, wboothprod1449, wboothprod1450, wadd1446d, wadd1446c );
smul_booth_prod u953 ( x[25], x[26], x[27], y[14], y[15], wboothprod1453 );
smul_booth_prod u954 ( x[27], x[28], x[29], y[12], y[13], wboothprod1454 );
smul_booth_prod u955 ( x[29], x[30], x[31], y[10], y[11], wboothprod1455 );
smul_full_add u956 ( wboothprod1453, wboothprod1454, wboothprod1455, wadd1451d, wadd1451c );
smul_half_add u957 ( wadd1446d, wadd1451d, wadd1444d, wadd1444c );
smul_full_add u958 ( wadd1431d, wadd1433d, wadd1444d, wadd1429d, wadd1429c );
smul_full_add u959 ( wadd1377c, wadd1425d, wadd1429d, wadd1423d, wadd1423c );
smul_half_add u960 ( wadd1375c, wadd1423d, wadd1421d, wadd1421c );
smul_carry_prop u961 ( wadd1332c, wadd1373d, wcarry1457g, wcarry1457p );
smul_carry_eval u962 ( wcarry1457g, wcarry1457p, wcarry1410, wcarry1456 );
smul_full_add u963 ( wadd1373c, wadd1421d, wcarry1456, wadd1419d, wadd1419c );
smul_full_add u964 ( wadd1431c, wadd1433c, wadd1444c, wadd1467d, wadd1467c );
smul_full_add u965 ( wadd1427c, wadd1429c, wadd1467d, wadd1465d, wadd1465c );
smul_full_add u966 ( wadd1435c, wadd1439c, wadd1446c, wadd1471d, wadd1471c );
smul_booth_prod u967 ( x[9], x[10], x[11], y[31], y[31], wboothprod1478 );
smul_inverter u968 ( wboothprod1478, winv1477 );
smul_booth_prod u969 ( x[11], x[12], x[13], y[29], y[30], wboothprod1479 );
smul_booth_prod u970 ( x[13], x[14], x[15], y[27], y[28], wboothprod1480 );
smul_full_add u971 ( winv1477, wboothprod1479, wboothprod1480, wadd1475d, wadd1475c );
smul_booth_prod u972 ( x[15], x[16], x[17], y[25], y[26], wboothprod1483 );
smul_booth_prod u973 ( x[17], x[18], x[19], y[23], y[24], wboothprod1484 );
smul_booth_prod u974 ( x[19], x[20], x[21], y[21], y[22], wboothprod1485 );
smul_full_add u975 ( wboothprod1483, wboothprod1484, wboothprod1485, wadd1481d, wadd1481c );
smul_full_add u976 ( wadd1451c, wadd1475d, wadd1481d, wadd1473d, wadd1473c );
smul_booth_prod u977 ( x[21], x[22], x[23], y[19], y[20], wboothprod1490 );
smul_booth_prod u978 ( x[23], x[24], x[25], y[17], y[18], wboothprod1491 );
smul_booth_prod u979 ( x[25], x[26], x[27], y[15], y[16], wboothprod1492 );
smul_full_add u980 ( wboothprod1490, wboothprod1491, wboothprod1492, wadd1488d, wadd1488c );
smul_booth_prod u981 ( x[27], x[28], x[29], y[13], y[14], wboothprod1493 );
smul_booth_prod u982 ( x[29], x[30], x[31], y[11], y[12], wboothprod1494 );
smul_full_add u983 ( wadd1488d, wboothprod1493, wboothprod1494, wadd1486d, wadd1486c );
smul_full_add u984 ( wadd1471d, wadd1473d, wadd1486d, wadd1469d, wadd1469c );
smul_full_add u985 ( wadd1425c, wadd1465d, wadd1469d, wadd1463d, wadd1463c );
smul_half_add u986 ( wadd1423c, wadd1463d, wadd1461d, wadd1461c );
smul_carry_prop u987 ( wadd1373c, wadd1421d, wcarry1498g, wcarry1498p );
smul_carry_merge u988 ( wcarry1457g, wcarry1457p, wcarry1498g, wcarry1498p, wcarry1496g, wcarry1496p );
smul_carry_eval u989 ( wcarry1496g, wcarry1496p, wcarry1410, wcarry1495 );
smul_full_add u990 ( wadd1421c, wadd1461d, wcarry1495, wadd1459d, wadd1459c );
smul_full_add u991 ( wadd1471c, wadd1473c, wadd1486c, wadd1508d, wadd1508c );
smul_full_add u992 ( wadd1467c, wadd1469c, wadd1508d, wadd1506d, wadd1506c );
smul_full_add u993 ( wadd1475c, wadd1481c, wadd1488c, wadd1512d, wadd1512c );
smul_booth_prod u994 ( x[11], x[12], x[13], y[30], y[31], wboothprod1518 );
smul_booth_prod u995 ( x[13], x[14], x[15], y[28], y[29], wboothprod1519 );
smul_full_add u996 ( 1'b1, wboothprod1518, wboothprod1519, wadd1516d, wadd1516c );
smul_booth_prod u997 ( x[15], x[16], x[17], y[26], y[27], wboothprod1522 );
smul_booth_prod u998 ( x[17], x[18], x[19], y[24], y[25], wboothprod1523 );
smul_booth_prod u999 ( x[19], x[20], x[21], y[22], y[23], wboothprod1524 );
smul_full_add u1000 ( wboothprod1522, wboothprod1523, wboothprod1524, wadd1520d, wadd1520c );
smul_booth_prod u1001 ( x[21], x[22], x[23], y[20], y[21], wboothprod1527 );
smul_booth_prod u1002 ( x[23], x[24], x[25], y[18], y[19], wboothprod1528 );
smul_booth_prod u1003 ( x[25], x[26], x[27], y[16], y[17], wboothprod1529 );
smul_full_add u1004 ( wboothprod1527, wboothprod1528, wboothprod1529, wadd1525d, wadd1525c );
smul_full_add u1005 ( wadd1516d, wadd1520d, wadd1525d, wadd1514d, wadd1514c );
smul_booth_prod u1006 ( x[27], x[28], x[29], y[14], y[15], wboothprod1532 );
smul_booth_prod u1007 ( x[29], x[30], x[31], y[12], y[13], wboothprod1533 );
smul_half_add u1008 ( wboothprod1532, wboothprod1533, wadd1530d, wadd1530c );
smul_full_add u1009 ( wadd1512d, wadd1514d, wadd1530d, wadd1510d, wadd1510c );
smul_full_add u1010 ( wadd1465c, wadd1506d, wadd1510d, wadd1504d, wadd1504c );
smul_half_add u1011 ( wadd1463c, wadd1504d, wadd1502d, wadd1502c );
smul_carry_prop u1012 ( wadd1421c, wadd1461d, wcarry1535g, wcarry1535p );
smul_carry_eval u1013 ( wcarry1535g, wcarry1535p, wcarry1495, wcarry1534 );
smul_full_add u1014 ( wadd1461c, wadd1502d, wcarry1534, wadd1500d, wadd1500c );
smul_full_add u1015 ( wadd1512c, wadd1514c, wadd1530c, wadd1545d, wadd1545c );
smul_full_add u1016 ( wadd1508c, wadd1510c, wadd1545d, wadd1543d, wadd1543c );
smul_full_add u1017 ( wadd1516c, wadd1520c, wadd1525c, wadd1549d, wadd1549c );
smul_booth_prod u1018 ( x[11], x[12], x[13], y[31], y[31], wboothprod1556 );
smul_inverter u1019 ( wboothprod1556, winv1555 );
smul_booth_prod u1020 ( x[13], x[14], x[15], y[29], y[30], wboothprod1557 );
smul_booth_prod u1021 ( x[15], x[16], x[17], y[27], y[28], wboothprod1558 );
smul_full_add u1022 ( winv1555, wboothprod1557, wboothprod1558, wadd1553d, wadd1553c );
smul_booth_prod u1023 ( x[17], x[18], x[19], y[25], y[26], wboothprod1561 );
smul_booth_prod u1024 ( x[19], x[20], x[21], y[23], y[24], wboothprod1562 );
smul_booth_prod u1025 ( x[21], x[22], x[23], y[21], y[22], wboothprod1563 );
smul_full_add u1026 ( wboothprod1561, wboothprod1562, wboothprod1563, wadd1559d, wadd1559c );
smul_booth_prod u1027 ( x[23], x[24], x[25], y[19], y[20], wboothprod1566 );
smul_booth_prod u1028 ( x[25], x[26], x[27], y[17], y[18], wboothprod1567 );
smul_booth_prod u1029 ( x[27], x[28], x[29], y[15], y[16], wboothprod1568 );
smul_full_add u1030 ( wboothprod1566, wboothprod1567, wboothprod1568, wadd1564d, wadd1564c );
smul_full_add u1031 ( wadd1553d, wadd1559d, wadd1564d, wadd1551d, wadd1551c );
smul_booth_prod u1032 ( x[29], x[30], x[31], y[13], y[14], wboothprod1569 );
smul_full_add u1033 ( wadd1549d, wadd1551d, wboothprod1569, wadd1547d, wadd1547c );
smul_full_add u1034 ( wadd1506c, wadd1543d, wadd1547d, wadd1541d, wadd1541c );
smul_half_add u1035 ( wadd1504c, wadd1541d, wadd1539d, wadd1539c );
smul_carry_prop u1036 ( wadd1461c, wadd1502d, wcarry1575g, wcarry1575p );
smul_carry_merge u1037 ( wcarry1535g, wcarry1535p, wcarry1575g, wcarry1575p, wcarry1573g, wcarry1573p );
smul_carry_merge u1038 ( wcarry1496g, wcarry1496p, wcarry1573g, wcarry1573p, wcarry1571g, wcarry1571p );
smul_carry_eval u1039 ( wcarry1571g, wcarry1571p, wcarry1410, wcarry1570 );
smul_full_add u1040 ( wadd1502c, wadd1539d, wcarry1570, wadd1537d, wadd1537c );
smul_full_add u1041 ( wadd1553c, wadd1559c, wadd1564c, wadd1587d, wadd1587c );
smul_full_add u1042 ( wadd1549c, wadd1551c, wadd1587d, wadd1585d, wadd1585c );
smul_full_add u1043 ( wadd1545c, wadd1547c, wadd1585d, wadd1583d, wadd1583c );
smul_booth_prod u1044 ( x[13], x[14], x[15], y[30], y[31], wboothprod1595 );
smul_booth_prod u1045 ( x[15], x[16], x[17], y[28], y[29], wboothprod1596 );
smul_full_add u1046 ( 1'b1, wboothprod1595, wboothprod1596, wadd1593d, wadd1593c );
smul_booth_prod u1047 ( x[17], x[18], x[19], y[26], y[27], wboothprod1599 );
smul_booth_prod u1048 ( x[19], x[20], x[21], y[24], y[25], wboothprod1600 );
smul_booth_prod u1049 ( x[21], x[22], x[23], y[22], y[23], wboothprod1601 );
smul_full_add u1050 ( wboothprod1599, wboothprod1600, wboothprod1601, wadd1597d, wadd1597c );
smul_booth_prod u1051 ( x[23], x[24], x[25], y[20], y[21], wboothprod1604 );
smul_booth_prod u1052 ( x[25], x[26], x[27], y[18], y[19], wboothprod1605 );
smul_booth_prod u1053 ( x[27], x[28], x[29], y[16], y[17], wboothprod1606 );
smul_full_add u1054 ( wboothprod1604, wboothprod1605, wboothprod1606, wadd1602d, wadd1602c );
smul_full_add u1055 ( wadd1593d, wadd1597d, wadd1602d, wadd1591d, wadd1591c );
smul_booth_prod u1056 ( x[29], x[30], x[31], y[14], y[15], wboothprod1607 );
smul_half_add u1057 ( wadd1591d, wboothprod1607, wadd1589d, wadd1589c );
smul_full_add u1058 ( wadd1543c, wadd1583d, wadd1589d, wadd1581d, wadd1581c );
smul_half_add u1059 ( wadd1541c, wadd1581d, wadd1579d, wadd1579c );
smul_carry_prop u1060 ( wadd1502c, wadd1539d, wcarry1609g, wcarry1609p );
smul_carry_eval u1061 ( wcarry1609g, wcarry1609p, wcarry1570, wcarry1608 );
smul_full_add u1062 ( wadd1539c, wadd1579d, wcarry1608, wadd1577d, wadd1577c );
smul_full_add u1063 ( wadd1593c, wadd1597c, wadd1602c, wadd1621d, wadd1621c );
smul_full_add u1064 ( wadd1587c, wadd1591c, wadd1621d, wadd1619d, wadd1619c );
smul_booth_prod u1065 ( x[13], x[14], x[15], y[31], y[31], wboothprod1628 );
smul_inverter u1066 ( wboothprod1628, winv1627 );
smul_booth_prod u1067 ( x[15], x[16], x[17], y[29], y[30], wboothprod1629 );
smul_booth_prod u1068 ( x[17], x[18], x[19], y[27], y[28], wboothprod1630 );
smul_full_add u1069 ( winv1627, wboothprod1629, wboothprod1630, wadd1625d, wadd1625c );
smul_booth_prod u1070 ( x[19], x[20], x[21], y[25], y[26], wboothprod1633 );
smul_booth_prod u1071 ( x[21], x[22], x[23], y[23], y[24], wboothprod1634 );
smul_booth_prod u1072 ( x[23], x[24], x[25], y[21], y[22], wboothprod1635 );
smul_full_add u1073 ( wboothprod1633, wboothprod1634, wboothprod1635, wadd1631d, wadd1631c );
smul_booth_prod u1074 ( x[25], x[26], x[27], y[19], y[20], wboothprod1638 );
smul_booth_prod u1075 ( x[27], x[28], x[29], y[17], y[18], wboothprod1639 );
smul_booth_prod u1076 ( x[29], x[30], x[31], y[15], y[16], wboothprod1640 );
smul_full_add u1077 ( wboothprod1638, wboothprod1639, wboothprod1640, wadd1636d, wadd1636c );
smul_full_add u1078 ( wadd1625d, wadd1631d, wadd1636d, wadd1623d, wadd1623c );
smul_full_add u1079 ( wadd1585c, wadd1619d, wadd1623d, wadd1617d, wadd1617c );
smul_full_add u1080 ( wadd1583c, wadd1589c, wadd1617d, wadd1615d, wadd1615c );
smul_half_add u1081 ( wadd1581c, wadd1615d, wadd1613d, wadd1613c );
smul_carry_prop u1082 ( wadd1539c, wadd1579d, wcarry1644g, wcarry1644p );
smul_carry_merge u1083 ( wcarry1609g, wcarry1609p, wcarry1644g, wcarry1644p, wcarry1642g, wcarry1642p );
smul_carry_eval u1084 ( wcarry1642g, wcarry1642p, wcarry1570, wcarry1641 );
smul_full_add u1085 ( wadd1579c, wadd1613d, wcarry1641, wadd1611d, wadd1611c );
smul_full_add u1086 ( wadd1625c, wadd1631c, wadd1636c, wadd1654d, wadd1654c );
smul_full_add u1087 ( wadd1621c, wadd1623c, wadd1654d, wadd1652d, wadd1652c );
smul_booth_prod u1088 ( x[15], x[16], x[17], y[30], y[31], wboothprod1660 );
smul_booth_prod u1089 ( x[17], x[18], x[19], y[28], y[29], wboothprod1661 );
smul_full_add u1090 ( 1'b1, wboothprod1660, wboothprod1661, wadd1658d, wadd1658c );
smul_booth_prod u1091 ( x[19], x[20], x[21], y[26], y[27], wboothprod1664 );
smul_booth_prod u1092 ( x[21], x[22], x[23], y[24], y[25], wboothprod1665 );
smul_booth_prod u1093 ( x[23], x[24], x[25], y[22], y[23], wboothprod1666 );
smul_full_add u1094 ( wboothprod1664, wboothprod1665, wboothprod1666, wadd1662d, wadd1662c );
smul_booth_prod u1095 ( x[25], x[26], x[27], y[20], y[21], wboothprod1669 );
smul_booth_prod u1096 ( x[27], x[28], x[29], y[18], y[19], wboothprod1670 );
smul_booth_prod u1097 ( x[29], x[30], x[31], y[16], y[17], wboothprod1671 );
smul_full_add u1098 ( wboothprod1669, wboothprod1670, wboothprod1671, wadd1667d, wadd1667c );
smul_full_add u1099 ( wadd1658d, wadd1662d, wadd1667d, wadd1656d, wadd1656c );
smul_full_add u1100 ( wadd1619c, wadd1652d, wadd1656d, wadd1650d, wadd1650c );
smul_full_add u1101 ( wadd1615c, wadd1617c, wadd1650d, wadd1648d, wadd1648c );
smul_carry_prop u1102 ( wadd1579c, wadd1613d, wcarry1673g, wcarry1673p );
smul_carry_eval u1103 ( wcarry1673g, wcarry1673p, wcarry1641, wcarry1672 );
smul_full_add u1104 ( wadd1613c, wadd1648d, wcarry1672, wadd1646d, wadd1646c );
smul_full_add u1105 ( wadd1658c, wadd1662c, wadd1667c, wadd1683d, wadd1683c );
smul_full_add u1106 ( wadd1654c, wadd1656c, wadd1683d, wadd1681d, wadd1681c );
smul_booth_prod u1107 ( x[15], x[16], x[17], y[31], y[31], wboothprod1690 );
smul_inverter u1108 ( wboothprod1690, winv1689 );
smul_booth_prod u1109 ( x[17], x[18], x[19], y[29], y[30], wboothprod1691 );
smul_booth_prod u1110 ( x[19], x[20], x[21], y[27], y[28], wboothprod1692 );
smul_full_add u1111 ( winv1689, wboothprod1691, wboothprod1692, wadd1687d, wadd1687c );
smul_booth_prod u1112 ( x[21], x[22], x[23], y[25], y[26], wboothprod1695 );
smul_booth_prod u1113 ( x[23], x[24], x[25], y[23], y[24], wboothprod1696 );
smul_booth_prod u1114 ( x[25], x[26], x[27], y[21], y[22], wboothprod1697 );
smul_full_add u1115 ( wboothprod1695, wboothprod1696, wboothprod1697, wadd1693d, wadd1693c );
smul_booth_prod u1116 ( x[27], x[28], x[29], y[19], y[20], wboothprod1700 );
smul_booth_prod u1117 ( x[29], x[30], x[31], y[17], y[18], wboothprod1701 );
smul_half_add u1118 ( wboothprod1700, wboothprod1701, wadd1698d, wadd1698c );
smul_full_add u1119 ( wadd1687d, wadd1693d, wadd1698d, wadd1685d, wadd1685c );
smul_full_add u1120 ( wadd1652c, wadd1681d, wadd1685d, wadd1679d, wadd1679c );
smul_half_add u1121 ( wadd1650c, wadd1679d, wadd1677d, wadd1677c );
smul_carry_prop u1122 ( wadd1613c, wadd1648d, wcarry1711g, wcarry1711p );
smul_carry_merge u1123 ( wcarry1673g, wcarry1673p, wcarry1711g, wcarry1711p, wcarry1709g, wcarry1709p );
smul_carry_merge u1124 ( wcarry1642g, wcarry1642p, wcarry1709g, wcarry1709p, wcarry1707g, wcarry1707p );
smul_carry_merge u1125 ( wcarry1571g, wcarry1571p, wcarry1707g, wcarry1707p, wcarry1705g, wcarry1705p );
smul_carry_merge u1126 ( wcarry1411g, wcarry1411p, wcarry1705g, wcarry1705p, wcarry1703g, wcarry1703p );
smul_carry_eval u1127 ( wcarry1703g, wcarry1703p, wcarry1025, wcarry1702 );
smul_full_add u1128 ( wadd1648c, wadd1677d, wcarry1702, wadd1675d, wadd1675c );
smul_full_add u1129 ( wadd1687c, wadd1693c, wadd1698c, wadd1721d, wadd1721c );
smul_full_add u1130 ( wadd1683c, wadd1685c, wadd1721d, wadd1719d, wadd1719c );
smul_booth_prod u1131 ( x[17], x[18], x[19], y[30], y[31], wboothprod1727 );
smul_booth_prod u1132 ( x[19], x[20], x[21], y[28], y[29], wboothprod1728 );
smul_full_add u1133 ( 1'b1, wboothprod1727, wboothprod1728, wadd1725d, wadd1725c );
smul_booth_prod u1134 ( x[21], x[22], x[23], y[26], y[27], wboothprod1731 );
smul_booth_prod u1135 ( x[23], x[24], x[25], y[24], y[25], wboothprod1732 );
smul_booth_prod u1136 ( x[25], x[26], x[27], y[22], y[23], wboothprod1733 );
smul_full_add u1137 ( wboothprod1731, wboothprod1732, wboothprod1733, wadd1729d, wadd1729c );
smul_booth_prod u1138 ( x[27], x[28], x[29], y[20], y[21], wboothprod1736 );
smul_booth_prod u1139 ( x[29], x[30], x[31], y[18], y[19], wboothprod1737 );
smul_half_add u1140 ( wboothprod1736, wboothprod1737, wadd1734d, wadd1734c );
smul_full_add u1141 ( wadd1725d, wadd1729d, wadd1734d, wadd1723d, wadd1723c );
smul_full_add u1142 ( wadd1681c, wadd1719d, wadd1723d, wadd1717d, wadd1717c );
smul_half_add u1143 ( wadd1679c, wadd1717d, wadd1715d, wadd1715c );
smul_carry_prop u1144 ( wadd1648c, wadd1677d, wcarry1739g, wcarry1739p );
smul_carry_eval u1145 ( wcarry1739g, wcarry1739p, wcarry1702, wcarry1738 );
smul_full_add u1146 ( wadd1677c, wadd1715d, wcarry1738, wadd1713d, wadd1713c );
smul_full_add u1147 ( wadd1725c, wadd1729c, wadd1734c, wadd1749d, wadd1749c );
smul_full_add u1148 ( wadd1721c, wadd1723c, wadd1749d, wadd1747d, wadd1747c );
smul_booth_prod u1149 ( x[17], x[18], x[19], y[31], y[31], wboothprod1756 );
smul_inverter u1150 ( wboothprod1756, winv1755 );
smul_booth_prod u1151 ( x[19], x[20], x[21], y[29], y[30], wboothprod1757 );
smul_booth_prod u1152 ( x[21], x[22], x[23], y[27], y[28], wboothprod1758 );
smul_full_add u1153 ( winv1755, wboothprod1757, wboothprod1758, wadd1753d, wadd1753c );
smul_booth_prod u1154 ( x[23], x[24], x[25], y[25], y[26], wboothprod1761 );
smul_booth_prod u1155 ( x[25], x[26], x[27], y[23], y[24], wboothprod1762 );
smul_booth_prod u1156 ( x[27], x[28], x[29], y[21], y[22], wboothprod1763 );
smul_full_add u1157 ( wboothprod1761, wboothprod1762, wboothprod1763, wadd1759d, wadd1759c );
smul_booth_prod u1158 ( x[29], x[30], x[31], y[19], y[20], wboothprod1764 );
smul_full_add u1159 ( wadd1753d, wadd1759d, wboothprod1764, wadd1751d, wadd1751c );
smul_full_add u1160 ( wadd1719c, wadd1747d, wadd1751d, wadd1745d, wadd1745c );
smul_half_add u1161 ( wadd1717c, wadd1745d, wadd1743d, wadd1743c );
smul_carry_prop u1162 ( wadd1677c, wadd1715d, wcarry1768g, wcarry1768p );
smul_carry_merge u1163 ( wcarry1739g, wcarry1739p, wcarry1768g, wcarry1768p, wcarry1766g, wcarry1766p );
smul_carry_eval u1164 ( wcarry1766g, wcarry1766p, wcarry1702, wcarry1765 );
smul_full_add u1165 ( wadd1715c, wadd1743d, wcarry1765, wadd1741d, wadd1741c );
smul_booth_prod u1166 ( x[19], x[20], x[21], y[30], y[31], wboothprod1782 );
smul_booth_prod u1167 ( x[21], x[22], x[23], y[28], y[29], wboothprod1783 );
smul_full_add u1168 ( 1'b1, wboothprod1782, wboothprod1783, wadd1780d, wadd1780c );
smul_full_add u1169 ( wadd1753c, wadd1759c, wadd1780d, wadd1778d, wadd1778c );
smul_full_add u1170 ( wadd1749c, wadd1751c, wadd1778d, wadd1776d, wadd1776c );
smul_booth_prod u1171 ( x[23], x[24], x[25], y[26], y[27], wboothprod1788 );
smul_booth_prod u1172 ( x[25], x[26], x[27], y[24], y[25], wboothprod1789 );
smul_booth_prod u1173 ( x[27], x[28], x[29], y[22], y[23], wboothprod1790 );
smul_full_add u1174 ( wboothprod1788, wboothprod1789, wboothprod1790, wadd1786d, wadd1786c );
smul_booth_prod u1175 ( x[29], x[30], x[31], y[20], y[21], wboothprod1791 );
smul_half_add u1176 ( wadd1786d, wboothprod1791, wadd1784d, wadd1784c );
smul_full_add u1177 ( wadd1747c, wadd1776d, wadd1784d, wadd1774d, wadd1774c );
smul_half_add u1178 ( wadd1745c, wadd1774d, wadd1772d, wadd1772c );
smul_carry_prop u1179 ( wadd1715c, wadd1743d, wcarry1793g, wcarry1793p );
smul_carry_eval u1180 ( wcarry1793g, wcarry1793p, wcarry1765, wcarry1792 );
smul_full_add u1181 ( wadd1743c, wadd1772d, wcarry1792, wadd1770d, wadd1770c );
smul_booth_prod u1182 ( x[19], x[20], x[21], y[31], y[31], wboothprod1808 );
smul_inverter u1183 ( wboothprod1808, winv1807 );
smul_booth_prod u1184 ( x[21], x[22], x[23], y[29], y[30], wboothprod1809 );
smul_booth_prod u1185 ( x[23], x[24], x[25], y[27], y[28], wboothprod1810 );
smul_full_add u1186 ( winv1807, wboothprod1809, wboothprod1810, wadd1805d, wadd1805c );
smul_full_add u1187 ( wadd1780c, wadd1786c, wadd1805d, wadd1803d, wadd1803c );
smul_booth_prod u1188 ( x[25], x[26], x[27], y[25], y[26], wboothprod1813 );
smul_booth_prod u1189 ( x[27], x[28], x[29], y[23], y[24], wboothprod1814 );
smul_booth_prod u1190 ( x[29], x[30], x[31], y[21], y[22], wboothprod1815 );
smul_full_add u1191 ( wboothprod1813, wboothprod1814, wboothprod1815, wadd1811d, wadd1811c );
smul_full_add u1192 ( wadd1778c, wadd1803d, wadd1811d, wadd1801d, wadd1801c );
smul_full_add u1193 ( wadd1776c, wadd1784c, wadd1801d, wadd1799d, wadd1799c );
smul_half_add u1194 ( wadd1774c, wadd1799d, wadd1797d, wadd1797c );
smul_carry_prop u1195 ( wadd1743c, wadd1772d, wcarry1821g, wcarry1821p );
smul_carry_merge u1196 ( wcarry1793g, wcarry1793p, wcarry1821g, wcarry1821p, wcarry1819g, wcarry1819p );
smul_carry_merge u1197 ( wcarry1766g, wcarry1766p, wcarry1819g, wcarry1819p, wcarry1817g, wcarry1817p );
smul_carry_eval u1198 ( wcarry1817g, wcarry1817p, wcarry1702, wcarry1816 );
smul_full_add u1199 ( wadd1772c, wadd1797d, wcarry1816, wadd1795d, wadd1795c );
smul_booth_prod u1200 ( x[21], x[22], x[23], y[30], y[31], wboothprod1833 );
smul_booth_prod u1201 ( x[23], x[24], x[25], y[28], y[29], wboothprod1834 );
smul_full_add u1202 ( 1'b1, wboothprod1833, wboothprod1834, wadd1831d, wadd1831c );
smul_full_add u1203 ( wadd1805c, wadd1811c, wadd1831d, wadd1829d, wadd1829c );
smul_booth_prod u1204 ( x[25], x[26], x[27], y[26], y[27], wboothprod1837 );
smul_booth_prod u1205 ( x[27], x[28], x[29], y[24], y[25], wboothprod1838 );
smul_booth_prod u1206 ( x[29], x[30], x[31], y[22], y[23], wboothprod1839 );
smul_full_add u1207 ( wboothprod1837, wboothprod1838, wboothprod1839, wadd1835d, wadd1835c );
smul_full_add u1208 ( wadd1803c, wadd1829d, wadd1835d, wadd1827d, wadd1827c );
smul_full_add u1209 ( wadd1799c, wadd1801c, wadd1827d, wadd1825d, wadd1825c );
smul_carry_prop u1210 ( wadd1772c, wadd1797d, wcarry1841g, wcarry1841p );
smul_carry_eval u1211 ( wcarry1841g, wcarry1841p, wcarry1816, wcarry1840 );
smul_full_add u1212 ( wadd1797c, wadd1825d, wcarry1840, wadd1823d, wadd1823c );
smul_booth_prod u1213 ( x[21], x[22], x[23], y[31], y[31], wboothprod1854 );
smul_inverter u1214 ( wboothprod1854, winv1853 );
smul_booth_prod u1215 ( x[23], x[24], x[25], y[29], y[30], wboothprod1855 );
smul_booth_prod u1216 ( x[25], x[26], x[27], y[27], y[28], wboothprod1856 );
smul_full_add u1217 ( winv1853, wboothprod1855, wboothprod1856, wadd1851d, wadd1851c );
smul_full_add u1218 ( wadd1831c, wadd1835c, wadd1851d, wadd1849d, wadd1849c );
smul_booth_prod u1219 ( x[27], x[28], x[29], y[25], y[26], wboothprod1859 );
smul_booth_prod u1220 ( x[29], x[30], x[31], y[23], y[24], wboothprod1860 );
smul_half_add u1221 ( wboothprod1859, wboothprod1860, wadd1857d, wadd1857c );
smul_full_add u1222 ( wadd1829c, wadd1849d, wadd1857d, wadd1847d, wadd1847c );
smul_full_add u1223 ( wadd1825c, wadd1827c, wadd1847d, wadd1845d, wadd1845c );
smul_carry_prop u1224 ( wadd1797c, wadd1825d, wcarry1864g, wcarry1864p );
smul_carry_merge u1225 ( wcarry1841g, wcarry1841p, wcarry1864g, wcarry1864p, wcarry1862g, wcarry1862p );
smul_carry_eval u1226 ( wcarry1862g, wcarry1862p, wcarry1816, wcarry1861 );
smul_full_add u1227 ( wadd1845d, 1'b0, wcarry1861, wadd1843d, wadd1843c );
smul_booth_prod u1228 ( x[23], x[24], x[25], y[30], y[31], wboothprod1876 );
smul_booth_prod u1229 ( x[25], x[26], x[27], y[28], y[29], wboothprod1877 );
smul_full_add u1230 ( 1'b1, wboothprod1876, wboothprod1877, wadd1874d, wadd1874c );
smul_booth_prod u1231 ( x[27], x[28], x[29], y[26], y[27], wboothprod1880 );
smul_booth_prod u1232 ( x[29], x[30], x[31], y[24], y[25], wboothprod1881 );
smul_half_add u1233 ( wboothprod1880, wboothprod1881, wadd1878d, wadd1878c );
smul_full_add u1234 ( wadd1851c, wadd1874d, wadd1878d, wadd1872d, wadd1872c );
smul_full_add u1235 ( wadd1849c, wadd1857c, wadd1872d, wadd1870d, wadd1870c );
smul_half_add u1236 ( wadd1847c, wadd1870d, wadd1868d, wadd1868c );
smul_carry_prop u1237 ( wadd1845d, 1'b0, wcarry1883g, wcarry1883p );
smul_carry_eval u1238 ( wcarry1883g, wcarry1883p, wcarry1861, wcarry1882 );
smul_full_add u1239 ( wadd1845c, wadd1868d, wcarry1882, wadd1866d, wadd1866c );
smul_booth_prod u1240 ( x[23], x[24], x[25], y[31], y[31], wboothprod1896 );
smul_inverter u1241 ( wboothprod1896, winv1895 );
smul_booth_prod u1242 ( x[25], x[26], x[27], y[29], y[30], wboothprod1897 );
smul_booth_prod u1243 ( x[27], x[28], x[29], y[27], y[28], wboothprod1898 );
smul_full_add u1244 ( winv1895, wboothprod1897, wboothprod1898, wadd1893d, wadd1893c );
smul_full_add u1245 ( wadd1874c, wadd1878c, wadd1893d, wadd1891d, wadd1891c );
smul_booth_prod u1246 ( x[29], x[30], x[31], y[25], y[26], wboothprod1899 );
smul_full_add u1247 ( wadd1872c, wadd1891d, wboothprod1899, wadd1889d, wadd1889c );
smul_half_add u1248 ( wadd1870c, wadd1889d, wadd1887d, wadd1887c );
smul_carry_prop u1249 ( wadd1845c, wadd1868d, wcarry1907g, wcarry1907p );
smul_carry_merge u1250 ( wcarry1883g, wcarry1883p, wcarry1907g, wcarry1907p, wcarry1905g, wcarry1905p );
smul_carry_merge u1251 ( wcarry1862g, wcarry1862p, wcarry1905g, wcarry1905p, wcarry1903g, wcarry1903p );
smul_carry_merge u1252 ( wcarry1817g, wcarry1817p, wcarry1903g, wcarry1903p, wcarry1901g, wcarry1901p );
smul_carry_eval u1253 ( wcarry1901g, wcarry1901p, wcarry1702, wcarry1900 );
smul_full_add u1254 ( wadd1868c, wadd1887d, wcarry1900, wadd1885d, wadd1885c );
smul_booth_prod u1255 ( x[25], x[26], x[27], y[30], y[31], wboothprod1917 );
smul_booth_prod u1256 ( x[27], x[28], x[29], y[28], y[29], wboothprod1918 );
smul_full_add u1257 ( 1'b1, wboothprod1917, wboothprod1918, wadd1915d, wadd1915c );
smul_booth_prod u1258 ( x[29], x[30], x[31], y[26], y[27], wboothprod1919 );
smul_full_add u1259 ( wadd1893c, wadd1915d, wboothprod1919, wadd1913d, wadd1913c );
smul_full_add u1260 ( wadd1889c, wadd1891c, wadd1913d, wadd1911d, wadd1911c );
smul_carry_prop u1261 ( wadd1868c, wadd1887d, wcarry1921g, wcarry1921p );
smul_carry_eval u1262 ( wcarry1921g, wcarry1921p, wcarry1900, wcarry1920 );
smul_full_add u1263 ( wadd1887c, wadd1911d, wcarry1920, wadd1909d, wadd1909c );
smul_booth_prod u1264 ( x[25], x[26], x[27], y[31], y[31], wboothprod1930 );
smul_inverter u1265 ( wboothprod1930, winv1929 );
smul_booth_prod u1266 ( x[27], x[28], x[29], y[29], y[30], wboothprod1931 );
smul_booth_prod u1267 ( x[29], x[30], x[31], y[27], y[28], wboothprod1932 );
smul_full_add u1268 ( winv1929, wboothprod1931, wboothprod1932, wadd1927d, wadd1927c );
smul_full_add u1269 ( wadd1913c, wadd1915c, wadd1927d, wadd1925d, wadd1925c );
smul_carry_prop u1270 ( wadd1887c, wadd1911d, wcarry1936g, wcarry1936p );
smul_carry_merge u1271 ( wcarry1921g, wcarry1921p, wcarry1936g, wcarry1936p, wcarry1934g, wcarry1934p );
smul_carry_eval u1272 ( wcarry1934g, wcarry1934p, wcarry1900, wcarry1933 );
smul_full_add u1273 ( wadd1911c, wadd1925d, wcarry1933, wadd1923d, wadd1923c );
smul_booth_prod u1274 ( x[27], x[28], x[29], y[30], y[31], wboothprod1944 );
smul_booth_prod u1275 ( x[29], x[30], x[31], y[28], y[29], wboothprod1945 );
smul_full_add u1276 ( 1'b1, wboothprod1944, wboothprod1945, wadd1942d, wadd1942c );
smul_full_add u1277 ( wadd1925c, wadd1927c, wadd1942d, wadd1940d, wadd1940c );
smul_carry_prop u1278 ( wadd1911c, wadd1925d, wcarry1947g, wcarry1947p );
smul_carry_eval u1279 ( wcarry1947g, wcarry1947p, wcarry1933, wcarry1946 );
smul_full_add u1280 ( wadd1940d, 1'b0, wcarry1946, wadd1938d, wadd1938c );
smul_booth_prod u1281 ( x[27], x[28], x[29], y[31], y[31], wboothprod1954 );
smul_inverter u1282 ( wboothprod1954, winv1953 );
smul_booth_prod u1283 ( x[29], x[30], x[31], y[29], y[30], wboothprod1955 );
smul_full_add u1284 ( wadd1942c, winv1953, wboothprod1955, wadd1951d, wadd1951c );
smul_carry_prop u1285 ( wadd1940d, 1'b0, wcarry1961g, wcarry1961p );
smul_carry_merge u1286 ( wcarry1947g, wcarry1947p, wcarry1961g, wcarry1961p, wcarry1959g, wcarry1959p );
smul_carry_merge u1287 ( wcarry1934g, wcarry1934p, wcarry1959g, wcarry1959p, wcarry1957g, wcarry1957p );
smul_carry_eval u1288 ( wcarry1957g, wcarry1957p, wcarry1900, wcarry1956 );
smul_full_add u1289 ( wadd1940c, wadd1951d, wcarry1956, wadd1949d, wadd1949c );
smul_booth_prod u1290 ( x[29], x[30], x[31], y[30], y[31], wboothprod1967 );
smul_full_add u1291 ( wadd1951c, 1'b1, wboothprod1967, wadd1965d, wadd1965c );
smul_carry_prop u1292 ( wadd1940c, wadd1951d, wcarry1969g, wcarry1969p );
smul_carry_eval u1293 ( wcarry1969g, wcarry1969p, wcarry1956, wcarry1968 );
smul_full_add u1294 ( wadd1965d, 1'b0, wcarry1968, wadd1963d, wadd1963c );
smul_booth_prod u1295 ( x[29], x[30], x[31], y[31], y[31], wboothprod1974 );
smul_inverter u1296 ( wboothprod1974, winv1973 );
smul_carry_prop u1297 ( wadd1965d, 1'b0, wcarry1978g, wcarry1978p );
smul_carry_merge u1298 ( wcarry1969g, wcarry1969p, wcarry1978g, wcarry1978p, wcarry1976g, wcarry1976p );
smul_carry_eval u1299 ( wcarry1976g, wcarry1976p, wcarry1956, wcarry1975 );
smul_full_add u1300 ( wadd1965c, winv1973, wcarry1975, wadd1971d, wadd1971c );
smul_carry_prop u1301 ( wadd1965c, winv1973, wcarry1983g, wcarry1983p );
smul_carry_eval u1302 ( wcarry1983g, wcarry1983p, wcarry1975, wcarry1982 );
smul_full_add u1303 ( 1'b1, 1'b0, wcarry1982, wadd1980d, wadd1980c );

assign p[0] = wadd0d;
assign p[1] = wadd4d;
assign p[2] = wadd10d;
assign p[3] = wadd22d;
assign p[4] = wadd31d;
assign p[5] = wadd48d;
assign p[6] = wadd60d;
assign p[7] = wadd78d;
assign p[8] = wadd93d;
assign p[9] = wadd118d;
assign p[10] = wadd136d;
assign p[11] = wadd160d;
assign p[12] = wadd181d;
assign p[13] = wadd210d;
assign p[14] = wadd234d;
assign p[15] = wadd264d;
assign p[16] = wadd291d;
assign p[17] = wadd330d;
assign p[18] = wadd360d;
assign p[19] = wadd396d;
assign p[20] = wadd429d;
assign p[21] = wadd470d;
assign p[22] = wadd506d;
assign p[23] = wadd548d;
assign p[24] = wadd587d;
assign p[25] = wadd636d;
assign p[26] = wadd678d;
assign p[27] = wadd726d;
assign p[28] = wadd771d;
assign p[29] = wadd824d;
assign p[30] = wadd872d;
assign p[31] = wadd926d;
assign p[32] = wadd977d;
assign p[33] = wadd1038d;
assign p[34] = wadd1088d;
assign p[35] = wadd1142d;
assign p[36] = wadd1189d;
assign p[37] = wadd1239d;
assign p[38] = wadd1283d;
assign p[39] = wadd1330d;
assign p[40] = wadd1371d;
assign p[41] = wadd1419d;
assign p[42] = wadd1459d;
assign p[43] = wadd1500d;
assign p[44] = wadd1537d;
assign p[45] = wadd1577d;
assign p[46] = wadd1611d;
assign p[47] = wadd1646d;
assign p[48] = wadd1675d;
assign p[49] = wadd1713d;
assign p[50] = wadd1741d;
assign p[51] = wadd1770d;
assign p[52] = wadd1795d;
assign p[53] = wadd1823d;
assign p[54] = wadd1843d;
assign p[55] = wadd1866d;
assign p[56] = wadd1885d;
assign p[57] = wadd1909d;
assign p[58] = wadd1923d;
assign p[59] = wadd1938d;
assign p[60] = wadd1949d;
assign p[61] = wadd1963d;
assign p[62] = wadd1971d;
assign p[63] = wadd1980d;

endmodule
